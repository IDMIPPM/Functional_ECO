module top (out_0, out_1, out_2, out_3, out_4, out_5, out_6, out_7, out_8, out_9, out_10, new_out1, new_out2, new_out3, new_out4, new_out5, in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, in_17, in_18, in_19, in_20, in_21, in_22, in_23, in_24, in_25, in_26, in_27, in_28, in_29, in_30, in_31);
	input in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, in_17, in_18, in_19, in_20, in_21, in_22, in_23, in_24, in_25, in_26, in_27, in_28, in_29, in_30, in_31;
	output out_0, out_1, out_2, out_3, out_4, out_5, out_6, out_7, out_8, out_9, out_10, out_11, new_out1, new_out2, new_out3, new_out4, new_out5;
	wire gm_n100, gm_n1000, gm_n1001, gm_n1002, gm_n1003, gm_n1004, gm_n1005, gm_n1006, gm_n1007, gm_n1008, gm_n1009, gm_n101, gm_n1010, gm_n1011, gm_n1012, gm_n1013, gm_n1014, gm_n1015, gm_n1016, gm_n1017, gm_n1018, gm_n1019, gm_n102, gm_n1020, gm_n1021, gm_n1022, gm_n1023, gm_n1024, gm_n1025, gm_n1026, gm_n1027, gm_n1028, gm_n1029, gm_n103, gm_n1030, gm_n1031, gm_n1032, gm_n1033, gm_n1034, gm_n1035, gm_n1036, gm_n1037, gm_n1038, gm_n1039, gm_n104, gm_n1040, gm_n1041, gm_n1042, gm_n1043, gm_n1044, gm_n1045, gm_n1046, gm_n1047, gm_n1048, gm_n1049, gm_n105, gm_n1050, gm_n1051, gm_n1052, gm_n1053, gm_n1054, gm_n1055, gm_n1056, gm_n1057, gm_n1058, gm_n1059, gm_n106, gm_n1060, gm_n1061, gm_n1062, gm_n1063, gm_n1064, gm_n1065, gm_n1066, gm_n1067, gm_n1068, gm_n1069, gm_n107, gm_n1070, gm_n1071, gm_n1072, gm_n1073, gm_n1074, gm_n1075, gm_n1076, gm_n1077, gm_n1078, gm_n1079, gm_n108, gm_n1080, gm_n1081, gm_n1082, gm_n1083, gm_n1084, gm_n1085, gm_n1086, gm_n1087, gm_n1088, gm_n1089, gm_n109, gm_n1090, gm_n1091, gm_n1092, gm_n1093, gm_n1094, gm_n1095, gm_n1096, gm_n1097, gm_n1098, gm_n1099, gm_n110, gm_n1100, gm_n1101, gm_n1102, gm_n1103, gm_n1104, gm_n1105, gm_n1106, gm_n1107, gm_n1108, gm_n1109, gm_n111, gm_n1110, gm_n1111, gm_n1112, gm_n1113, gm_n1114, gm_n1115, gm_n1116, gm_n1117, gm_n1118, gm_n1119, gm_n112, gm_n1120, gm_n1121, gm_n1122, gm_n1123, gm_n1124, gm_n1125, gm_n1126, gm_n1127, gm_n1128, gm_n1129, gm_n113, gm_n1130, gm_n1131, gm_n1132, gm_n1133, gm_n1134, gm_n1135, gm_n1136, gm_n1137, gm_n1138, gm_n1139, gm_n114, gm_n1140, gm_n1141, gm_n1142, gm_n1143, gm_n1144, gm_n1145, gm_n1146, gm_n1147, gm_n1148, gm_n1149, gm_n115, gm_n1150, gm_n1151, gm_n1152, gm_n1153, gm_n1154, gm_n1155, gm_n1156, gm_n1157, gm_n1158, gm_n1159, gm_n116, gm_n1160, gm_n1161, gm_n1162, gm_n1163, gm_n1164, gm_n1165, gm_n1166, gm_n1167, gm_n1168, gm_n1169, gm_n117, gm_n1170, gm_n1171, gm_n1172, gm_n1173, gm_n1174, gm_n1175, gm_n1176, gm_n1177, gm_n1178, gm_n1179, gm_n118, gm_n1180, gm_n1181, gm_n1182, gm_n1183, gm_n1184, gm_n1185, gm_n1186, gm_n1187, gm_n1188, gm_n1189, gm_n119, gm_n1190, gm_n1191, gm_n1192, gm_n1193, gm_n1194, gm_n1195, gm_n1196, gm_n1197, gm_n1198, gm_n1199, gm_n120, gm_n1200, gm_n1201, gm_n1202, gm_n1203, gm_n1204, gm_n1206, gm_n1207, gm_n1208, gm_n1209, gm_n121, gm_n1210, gm_n1211, gm_n1212, gm_n1213, gm_n1214, gm_n1215, gm_n1216, gm_n1217, gm_n1218, gm_n1219, gm_n122, gm_n1220, gm_n1221, gm_n1222, gm_n1223, gm_n1224, gm_n1225, gm_n1226, gm_n1227, gm_n1228, gm_n1229, gm_n123, gm_n1230, gm_n1231, gm_n1232, gm_n1233, gm_n1234, gm_n1235, gm_n1236, gm_n1237, gm_n1238, gm_n1239, gm_n124, gm_n1240, gm_n1241, gm_n1242, gm_n1243, gm_n1244, gm_n1245, gm_n1246, gm_n1247, gm_n1248, gm_n1249, gm_n125, gm_n1250, gm_n1251, gm_n1252, gm_n1253, gm_n1254, gm_n1255, gm_n1256, gm_n1257, gm_n1258, gm_n1259, gm_n126, gm_n1260, gm_n1261, gm_n1262, gm_n1263, gm_n1264, gm_n1265, gm_n1266, gm_n1267, gm_n1268, gm_n1269, gm_n127, gm_n1270, gm_n1271, gm_n1272, gm_n1273, gm_n1274, gm_n1275, gm_n1276, gm_n1277, gm_n1278, gm_n1279, gm_n128, gm_n1280, gm_n1281, gm_n1282, gm_n1283, gm_n1284, gm_n1285, gm_n1286, gm_n1287, gm_n1288, gm_n1289, gm_n129, gm_n1290, gm_n1291, gm_n1292, gm_n1293, gm_n1294, gm_n1295, gm_n1296, gm_n1297, gm_n1298, gm_n1299, gm_n130, gm_n1300, gm_n1301, gm_n1302, gm_n1303, gm_n1304, gm_n1305, gm_n1306, gm_n1307, gm_n1308, gm_n1309, gm_n131, gm_n1310, gm_n1311, gm_n1312, gm_n1313, gm_n1314, gm_n1315, gm_n1316, gm_n1317, gm_n1318, gm_n1319, gm_n132, gm_n1320, gm_n1321, gm_n1322, gm_n1323, gm_n1324, gm_n1325, gm_n1326, gm_n1327, gm_n1328, gm_n1329, gm_n133, gm_n1330, gm_n1331, gm_n1332, gm_n1333, gm_n1334, gm_n1335, gm_n1336, gm_n1337, gm_n1338, gm_n1339, gm_n134, gm_n1340, gm_n1341, gm_n1342, gm_n1343, gm_n1344, gm_n1345, gm_n1346, gm_n1347, gm_n1348, gm_n1349, gm_n135, gm_n1350, gm_n1351, gm_n1352, gm_n1353, gm_n1354, gm_n1355, gm_n1356, gm_n1357, gm_n1358, gm_n1359, gm_n136, gm_n1360, gm_n1361, gm_n1362, gm_n1363, gm_n1364, gm_n1365, gm_n1366, gm_n1367, gm_n1368, gm_n1369, gm_n137, gm_n1370, gm_n1371, gm_n1372, gm_n1373, gm_n1374, gm_n1375, gm_n1376, gm_n1377, gm_n1378, gm_n1379, gm_n138, gm_n1380, gm_n1381, gm_n1382, gm_n1383, gm_n1384, gm_n1385, gm_n1386, gm_n1387, gm_n1388, gm_n1389, gm_n139, gm_n1390, gm_n1391, gm_n1392, gm_n1393, gm_n1394, gm_n1395, gm_n1396, gm_n1397, gm_n1398, gm_n1399, gm_n140, gm_n1400, gm_n1401, gm_n1402, gm_n1403, gm_n1404, gm_n1405, gm_n1406, gm_n1407, gm_n1408, gm_n141, gm_n1410, gm_n1411, gm_n1412, gm_n1413, gm_n1414, gm_n1415, gm_n1416, gm_n1417, gm_n1418, gm_n1419, gm_n142, gm_n1420, gm_n1421, gm_n1422, gm_n1423, gm_n1424, gm_n1425, gm_n1426, gm_n1427, gm_n1428, gm_n1429, gm_n143, gm_n1430, gm_n1431, gm_n1432, gm_n1433, gm_n1434, gm_n1435, gm_n1436, gm_n1437, gm_n1438, gm_n1439, gm_n144, gm_n1440, gm_n1441, gm_n1442, gm_n1443, gm_n1444, gm_n1445, gm_n1446, gm_n1447, gm_n1448, gm_n1449, gm_n145, gm_n1450, gm_n1451, gm_n1452, gm_n1453, gm_n1454, gm_n1455, gm_n1456, gm_n1457, gm_n1458, gm_n1459, gm_n146, gm_n1460, gm_n1461, gm_n1462, gm_n1463, gm_n1464, gm_n1465, gm_n1466, gm_n1467, gm_n1468, gm_n1469, gm_n147, gm_n1470, gm_n1471, gm_n1472, gm_n1473, gm_n1474, gm_n1475, gm_n1476, gm_n1477, gm_n1478, gm_n1479, gm_n148, gm_n1480, gm_n1481, gm_n1482, gm_n1483, gm_n1484, gm_n1485, gm_n1486, gm_n1487, gm_n1488, gm_n1489, gm_n149, gm_n1490, gm_n1491, gm_n1492, gm_n1493, gm_n1494, gm_n1495, gm_n1496, gm_n1497, gm_n1498, gm_n1499, gm_n150, gm_n1500, gm_n1501, gm_n1502, gm_n1503, gm_n1504, gm_n1505, gm_n1506, gm_n1507, gm_n1508, gm_n1509, gm_n151, gm_n1510, gm_n1511, gm_n1512, gm_n1513, gm_n1514, gm_n1515, gm_n1516, gm_n1517, gm_n1518, gm_n1519, gm_n152, gm_n1520, gm_n1521, gm_n1522, gm_n1523, gm_n1524, gm_n1525, gm_n1526, gm_n1527, gm_n1528, gm_n1529, gm_n153, gm_n1530, gm_n1531, gm_n1532, gm_n1533, gm_n1534, gm_n1535, gm_n1536, gm_n1537, gm_n1538, gm_n1539, gm_n154, gm_n1540, gm_n1541, gm_n1542, gm_n1543, gm_n1544, gm_n1545, gm_n1546, gm_n1547, gm_n1548, gm_n1549, gm_n155, gm_n1550, gm_n1551, gm_n1552, gm_n1553, gm_n1554, gm_n1555, gm_n1556, gm_n1557, gm_n1558, gm_n1559, gm_n156, gm_n1560, gm_n1561, gm_n1562, gm_n1563, gm_n1564, gm_n1565, gm_n1566, gm_n1567, gm_n1568, gm_n1569, gm_n157, gm_n1570, gm_n1571, gm_n1572, gm_n1573, gm_n1574, gm_n1575, gm_n1576, gm_n1577, gm_n1578, gm_n1579, gm_n158, gm_n1580, gm_n1581, gm_n1582, gm_n1583, gm_n1584, gm_n1585, gm_n1586, gm_n1587, gm_n1588, gm_n1589, gm_n159, gm_n1590, gm_n1591, gm_n1592, gm_n1593, gm_n1594, gm_n1595, gm_n1596, gm_n1597, gm_n1598, gm_n1599, gm_n160, gm_n1600, gm_n1601, gm_n1602, gm_n1604, gm_n1605, gm_n1606, gm_n1607, gm_n1608, gm_n1609, gm_n161, gm_n1610, gm_n1611, gm_n1612, gm_n1613, gm_n1614, gm_n1615, gm_n1616, gm_n1617, gm_n1618, gm_n1619, gm_n162, gm_n1620, gm_n1621, gm_n1622, gm_n1623, gm_n1624, gm_n1625, gm_n1626, gm_n1627, gm_n1628, gm_n1629, gm_n163, gm_n1630, gm_n1631, gm_n1632, gm_n1633, gm_n1634, gm_n1635, gm_n1636, gm_n1637, gm_n1638, gm_n1639, gm_n164, gm_n1640, gm_n1641, gm_n1642, gm_n1643, gm_n1644, gm_n1645, gm_n1646, gm_n1647, gm_n1648, gm_n1649, gm_n165, gm_n1650, gm_n1651, gm_n1652, gm_n1653, gm_n1654, gm_n1655, gm_n1656, gm_n1657, gm_n1658, gm_n1659, gm_n166, gm_n1660, gm_n1661, gm_n1662, gm_n1663, gm_n1664, gm_n1665, gm_n1666, gm_n1667, gm_n1668, gm_n1669, gm_n167, gm_n1670, gm_n1671, gm_n1672, gm_n1673, gm_n1674, gm_n1675, gm_n1676, gm_n1677, gm_n1678, gm_n1679, gm_n168, gm_n1680, gm_n1681, gm_n1682, gm_n1683, gm_n1684, gm_n1685, gm_n1686, gm_n1687, gm_n1688, gm_n1689, gm_n169, gm_n1690, gm_n1691, gm_n1692, gm_n1693, gm_n1694, gm_n1695, gm_n1696, gm_n1697, gm_n1698, gm_n1699, gm_n170, gm_n1700, gm_n1701, gm_n1702, gm_n1703, gm_n1704, gm_n1705, gm_n1706, gm_n1707, gm_n1708, gm_n1709, gm_n171, gm_n1710, gm_n1711, gm_n1712, gm_n1713, gm_n1714, gm_n1715, gm_n1716, gm_n1717, gm_n1718, gm_n1719, gm_n172, gm_n1720, gm_n1721, gm_n1722, gm_n1723, gm_n1724, gm_n1725, gm_n1726, gm_n1727, gm_n1728, gm_n1729, gm_n173, gm_n1730, gm_n1731, gm_n1732, gm_n1733, gm_n1734, gm_n1735, gm_n1736, gm_n1737, gm_n1738, gm_n1739, gm_n174, gm_n1740, gm_n1741, gm_n1742, gm_n1743, gm_n1744, gm_n1745, gm_n1746, gm_n1747, gm_n1748, gm_n1749, gm_n175, gm_n1750, gm_n1751, gm_n1752, gm_n1753, gm_n1754, gm_n1755, gm_n1756, gm_n1757, gm_n1758, gm_n1759, gm_n176, gm_n1760, gm_n1761, gm_n1762, gm_n1763, gm_n1764, gm_n1765, gm_n1766, gm_n1767, gm_n1768, gm_n1769, gm_n177, gm_n1770, gm_n1771, gm_n1772, gm_n1773, gm_n1774, gm_n1775, gm_n1776, gm_n1777, gm_n1778, gm_n1779, gm_n178, gm_n1780, gm_n1781, gm_n1782, gm_n1783, gm_n1784, gm_n1785, gm_n1786, gm_n1787, gm_n1788, gm_n1789, gm_n179, gm_n1790, gm_n1791, gm_n1792, gm_n1793, gm_n1794, gm_n1795, gm_n1796, gm_n1797, gm_n1798, gm_n1799, gm_n180, gm_n1800, gm_n1801, gm_n1802, gm_n1803, gm_n1805, gm_n1806, gm_n1807, gm_n1808, gm_n1809, gm_n181, gm_n1810, gm_n1811, gm_n1812, gm_n1813, gm_n1814, gm_n1815, gm_n1816, gm_n1817, gm_n1818, gm_n1819, gm_n182, gm_n1820, gm_n1821, gm_n1822, gm_n1823, gm_n1824, gm_n1825, gm_n1826, gm_n1827, gm_n1828, gm_n1829, gm_n183, gm_n1830, gm_n1831, gm_n1832, gm_n1833, gm_n1834, gm_n1835, gm_n1836, gm_n1837, gm_n1838, gm_n1839, gm_n184, gm_n1840, gm_n1841, gm_n1842, gm_n1843, gm_n1844, gm_n1845, gm_n1846, gm_n1847, gm_n1848, gm_n1849, gm_n185, gm_n1850, gm_n1851, gm_n1852, gm_n1853, gm_n1854, gm_n1855, gm_n1856, gm_n1857, gm_n1858, gm_n1859, gm_n186, gm_n1860, gm_n1861, gm_n1862, gm_n1863, gm_n1864, gm_n1865, gm_n1866, gm_n1867, gm_n1868, gm_n1869, gm_n187, gm_n1870, gm_n1871, gm_n1872, gm_n1873, gm_n1874, gm_n1875, gm_n1876, gm_n1877, gm_n1878, gm_n1879, gm_n188, gm_n1880, gm_n1881, gm_n1882, gm_n1883, gm_n1884, gm_n1885, gm_n1886, gm_n1887, gm_n1888, gm_n1889, gm_n189, gm_n1890, gm_n1891, gm_n1892, gm_n1893, gm_n1894, gm_n1895, gm_n1896, gm_n1897, gm_n1898, gm_n1899, gm_n190, gm_n1900, gm_n1901, gm_n1902, gm_n1903, gm_n1904, gm_n1905, gm_n1906, gm_n1907, gm_n1908, gm_n1909, gm_n191, gm_n1910, gm_n1911, gm_n1912, gm_n1913, gm_n1914, gm_n1915, gm_n1916, gm_n1917, gm_n1918, gm_n1919, gm_n192, gm_n1920, gm_n1921, gm_n1922, gm_n1923, gm_n1924, gm_n1925, gm_n1926, gm_n1927, gm_n1928, gm_n1929, gm_n193, gm_n1930, gm_n1931, gm_n1932, gm_n1933, gm_n1934, gm_n1935, gm_n1936, gm_n1937, gm_n1938, gm_n1939, gm_n194, gm_n1940, gm_n1941, gm_n1942, gm_n1943, gm_n1944, gm_n1945, gm_n1946, gm_n1947, gm_n1948, gm_n1949, gm_n195, gm_n1950, gm_n1951, gm_n1952, gm_n1953, gm_n1954, gm_n1955, gm_n1956, gm_n1957, gm_n1958, gm_n1959, gm_n196, gm_n1960, gm_n1961, gm_n1962, gm_n1963, gm_n1964, gm_n1965, gm_n1966, gm_n1967, gm_n1968, gm_n1969, gm_n197, gm_n1970, gm_n1971, gm_n1972, gm_n1973, gm_n1974, gm_n1975, gm_n1976, gm_n1977, gm_n1978, gm_n1979, gm_n198, gm_n1980, gm_n1981, gm_n1982, gm_n1983, gm_n1984, gm_n1985, gm_n1986, gm_n1987, gm_n1988, gm_n1989, gm_n199, gm_n1990, gm_n1991, gm_n1992, gm_n1993, gm_n1994, gm_n1995, gm_n1996, gm_n1997, gm_n1998, gm_n1999, gm_n200, gm_n2000, gm_n2001, gm_n2002, gm_n2004, gm_n2005, gm_n2006, gm_n2007, gm_n2008, gm_n2009, gm_n201, gm_n2010, gm_n2011, gm_n2012, gm_n2013, gm_n2014, gm_n2015, gm_n2016, gm_n2017, gm_n2018, gm_n2019, gm_n202, gm_n2020, gm_n2021, gm_n2022, gm_n2023, gm_n2024, gm_n2025, gm_n2026, gm_n2027, gm_n2028, gm_n2029, gm_n203, gm_n2030, gm_n2031, gm_n2032, gm_n2033, gm_n2034, gm_n2035, gm_n2036, gm_n2037, gm_n2038, gm_n2039, gm_n204, gm_n2040, gm_n2041, gm_n2042, gm_n2043, gm_n2044, gm_n2045, gm_n2046, gm_n2047, gm_n2048, gm_n2049, gm_n205, gm_n2050, gm_n2051, gm_n2052, gm_n2053, gm_n2054, gm_n2055, gm_n2056, gm_n2057, gm_n2058, gm_n2059, gm_n206, gm_n2060, gm_n2061, gm_n2062, gm_n2063, gm_n2064, gm_n2065, gm_n2066, gm_n2067, gm_n2068, gm_n2069, gm_n207, gm_n2070, gm_n2071, gm_n2072, gm_n2073, gm_n2074, gm_n2075, gm_n2076, gm_n2077, gm_n2078, gm_n2079, gm_n208, gm_n2080, gm_n2081, gm_n2082, gm_n2083, gm_n2084, gm_n2085, gm_n2086, gm_n2087, gm_n2088, gm_n2089, gm_n209, gm_n2090, gm_n2091, gm_n2092, gm_n2093, gm_n2094, gm_n2095, gm_n2096, gm_n2097, gm_n2098, gm_n2099, gm_n210, gm_n2100, gm_n2101, gm_n2102, gm_n2103, gm_n2104, gm_n2105, gm_n2106, gm_n2107, gm_n2108, gm_n2109, gm_n211, gm_n2110, gm_n2111, gm_n2112, gm_n2113, gm_n2114, gm_n2115, gm_n2116, gm_n2117, gm_n2118, gm_n2119, gm_n212, gm_n2120, gm_n2121, gm_n2122, gm_n2123, gm_n2124, gm_n2125, gm_n2126, gm_n2127, gm_n2128, gm_n2129, gm_n213, gm_n2130, gm_n2131, gm_n2132, gm_n2133, gm_n2134, gm_n2135, gm_n2136, gm_n2137, gm_n2138, gm_n2139, gm_n214, gm_n2140, gm_n2141, gm_n2142, gm_n2143, gm_n2144, gm_n2145, gm_n2146, gm_n2147, gm_n2148, gm_n2149, gm_n215, gm_n2150, gm_n2151, gm_n2152, gm_n2153, gm_n2154, gm_n2155, gm_n2156, gm_n2157, gm_n2158, gm_n2159, gm_n216, gm_n2160, gm_n2161, gm_n2162, gm_n2163, gm_n2164, gm_n2165, gm_n2166, gm_n2167, gm_n2168, gm_n2169, gm_n217, gm_n2170, gm_n2171, gm_n2172, gm_n2173, gm_n2174, gm_n2175, gm_n2176, gm_n2177, gm_n2178, gm_n2179, gm_n218, gm_n2180, gm_n2181, gm_n2182, gm_n2183, gm_n2184, gm_n2185, gm_n2186, gm_n2187, gm_n2188, gm_n2189, gm_n219, gm_n2190, gm_n2191, gm_n2192, gm_n2193, gm_n2194, gm_n2195, gm_n2196, gm_n2198, gm_n2199, gm_n220, gm_n2200, gm_n2201, gm_n2202, gm_n2203, gm_n2204, gm_n2205, gm_n2206, gm_n2207, gm_n2208, gm_n2209, gm_n221, gm_n2210, gm_n2211, gm_n2212, gm_n2213, gm_n2214, gm_n2215, gm_n2216, gm_n2217, gm_n2218, gm_n2219, gm_n222, gm_n2220, gm_n2221, gm_n2222, gm_n2223, gm_n2224, gm_n2225, gm_n2226, gm_n2227, gm_n2228, gm_n2229, gm_n223, gm_n2230, gm_n2231, gm_n2232, gm_n2233, gm_n2234, gm_n2235, gm_n2236, gm_n2237, gm_n2238, gm_n2239, gm_n224, gm_n2240, gm_n2241, gm_n2242, gm_n2243, gm_n2244, gm_n2245, gm_n2246, gm_n2247, gm_n2248, gm_n2249, gm_n225, gm_n2250, gm_n2251, gm_n2252, gm_n2253, gm_n2254, gm_n2255, gm_n2256, gm_n2257, gm_n2258, gm_n2259, gm_n226, gm_n2260, gm_n2261, gm_n2262, gm_n2263, gm_n2264, gm_n2265, gm_n2266, gm_n2267, gm_n2268, gm_n2269, gm_n227, gm_n2270, gm_n2271, gm_n2272, gm_n2273, gm_n2274, gm_n2275, gm_n2276, gm_n2277, gm_n2278, gm_n2279, gm_n228, gm_n2280, gm_n2281, gm_n2282, gm_n2283, gm_n2284, gm_n2285, gm_n2286, gm_n2287, gm_n2288, gm_n2289, gm_n229, gm_n2290, gm_n2291, gm_n2292, gm_n2293, gm_n2294, gm_n2295, gm_n2296, gm_n2297, gm_n2298, gm_n2299, gm_n230, gm_n2300, gm_n2301, gm_n2302, gm_n2303, gm_n2304, gm_n2305, gm_n2306, gm_n2307, gm_n2308, gm_n2309, gm_n231, gm_n2310, gm_n2311, gm_n2312, gm_n2313, gm_n2314, gm_n2315, gm_n2316, gm_n2317, gm_n2318, gm_n2319, gm_n232, gm_n2320, gm_n2321, gm_n2322, gm_n2323, gm_n2324, gm_n2325, gm_n2326, gm_n2327, gm_n2328, gm_n2329, gm_n233, gm_n2330, gm_n2331, gm_n2332, gm_n2333, gm_n2334, gm_n2335, gm_n2336, gm_n2337, gm_n2338, gm_n2339, gm_n234, gm_n2340, gm_n2341, gm_n2342, gm_n2343, gm_n2344, gm_n2345, gm_n2346, gm_n2347, gm_n2348, gm_n2349, gm_n235, gm_n2350, gm_n2351, gm_n2352, gm_n2353, gm_n2354, gm_n2355, gm_n2356, gm_n2357, gm_n2358, gm_n2359, gm_n236, gm_n2360, gm_n2361, gm_n2362, gm_n2363, gm_n2364, gm_n2365, gm_n2366, gm_n2367, gm_n2368, gm_n2369, gm_n237, gm_n2370, gm_n2371, gm_n2372, gm_n2373, gm_n2374, gm_n2375, gm_n2376, gm_n2377, gm_n2378, gm_n2379, gm_n238, gm_n2381, gm_n2382, gm_n2383, gm_n2384, gm_n2385, gm_n2386, gm_n2387, gm_n2388, gm_n2389, gm_n239, gm_n2390, gm_n2391, gm_n2392, gm_n2393, gm_n2394, gm_n2395, gm_n2396, gm_n2397, gm_n2398, gm_n2399, gm_n240, gm_n2400, gm_n2401, gm_n2402, gm_n2403, gm_n2404, gm_n2405, gm_n2406, gm_n2407, gm_n2408, gm_n2409, gm_n241, gm_n2410, gm_n2411, gm_n2412, gm_n2413, gm_n2414, gm_n2415, gm_n2416, gm_n2417, gm_n2418, gm_n2419, gm_n242, gm_n2420, gm_n2421, gm_n2422, gm_n2423, gm_n2424, gm_n2425, gm_n2426, gm_n2427, gm_n2428, gm_n2429, gm_n243, gm_n2430, gm_n2431, gm_n2432, gm_n2433, gm_n2434, gm_n2435, gm_n2436, gm_n2437, gm_n2438, gm_n2439, gm_n244, gm_n2440, gm_n2441, gm_n2442, gm_n2443, gm_n2444, gm_n2445, gm_n2446, gm_n2447, gm_n2448, gm_n2449, gm_n245, gm_n2450, gm_n2451, gm_n2452, gm_n2453, gm_n2454, gm_n2455, gm_n2456, gm_n2457, gm_n2458, gm_n2459, gm_n246, gm_n2460, gm_n2461, gm_n2462, gm_n2463, gm_n2464, gm_n2465, gm_n2466, gm_n2467, gm_n2468, gm_n2469, gm_n247, gm_n2470, gm_n2471, gm_n2472, gm_n2473, gm_n2474, gm_n2475, gm_n2476, gm_n2477, gm_n2478, gm_n2479, gm_n248, gm_n2480, gm_n2481, gm_n2482, gm_n2483, gm_n2484, gm_n2485, gm_n2486, gm_n2487, gm_n2488, gm_n2489, gm_n249, gm_n2490, gm_n2491, gm_n2492, gm_n2493, gm_n2494, gm_n2495, gm_n2496, gm_n2497, gm_n2498, gm_n2499, gm_n250, gm_n2500, gm_n2501, gm_n2502, gm_n2503, gm_n2504, gm_n2505, gm_n2506, gm_n2507, gm_n2508, gm_n2509, gm_n251, gm_n2510, gm_n2511, gm_n2512, gm_n2513, gm_n2514, gm_n2515, gm_n2516, gm_n2517, gm_n2518, gm_n2519, gm_n252, gm_n2520, gm_n2521, gm_n2522, gm_n2523, gm_n2524, gm_n2525, gm_n2526, gm_n2527, gm_n2528, gm_n2529, gm_n253, gm_n2530, gm_n2531, gm_n2532, gm_n2533, gm_n2534, gm_n2535, gm_n2536, gm_n2537, gm_n2538, gm_n2539, gm_n254, gm_n2540, gm_n2541, gm_n2542, gm_n2543, gm_n2544, gm_n2545, gm_n2546, gm_n2547, gm_n2548, gm_n2549, gm_n255, gm_n2550, gm_n2551, gm_n2552, gm_n2553, gm_n2554, gm_n2555, gm_n2556, gm_n2557, gm_n2558, gm_n2559, gm_n256, gm_n2560, gm_n2561, gm_n2562, gm_n2564, gm_n2565, gm_n2566, gm_n2567, gm_n2568, gm_n2569, gm_n257, gm_n2570, gm_n2571, gm_n2572, gm_n2573, gm_n2574, gm_n2575, gm_n2576, gm_n2577, gm_n2578, gm_n2579, gm_n258, gm_n2580, gm_n2581, gm_n2582, gm_n2583, gm_n2584, gm_n2585, gm_n2586, gm_n2587, gm_n2588, gm_n2589, gm_n259, gm_n2590, gm_n2591, gm_n2592, gm_n2593, gm_n2594, gm_n2595, gm_n2596, gm_n2597, gm_n2598, gm_n2599, gm_n260, gm_n2600, gm_n2601, gm_n2602, gm_n2603, gm_n2604, gm_n2605, gm_n2606, gm_n2607, gm_n2608, gm_n2609, gm_n261, gm_n2610, gm_n2611, gm_n2612, gm_n2613, gm_n2614, gm_n2615, gm_n2616, gm_n2617, gm_n2618, gm_n2619, gm_n262, gm_n2620, gm_n2621, gm_n2622, gm_n2623, gm_n2624, gm_n2625, gm_n2626, gm_n2627, gm_n2628, gm_n2629, gm_n263, gm_n2630, gm_n2631, gm_n2632, gm_n2633, gm_n2634, gm_n2635, gm_n2636, gm_n2637, gm_n2638, gm_n2639, gm_n264, gm_n2640, gm_n2641, gm_n2642, gm_n2643, gm_n2644, gm_n2645, gm_n2646, gm_n2647, gm_n2648, gm_n2649, gm_n265, gm_n2650, gm_n2651, gm_n2652, gm_n2653, gm_n2654, gm_n2655, gm_n2656, gm_n2657, gm_n2658, gm_n2659, gm_n266, gm_n2660, gm_n2661, gm_n2662, gm_n2663, gm_n2664, gm_n2665, gm_n2666, gm_n2667, gm_n2668, gm_n2669, gm_n267, gm_n2670, gm_n2671, gm_n2672, gm_n2673, gm_n2674, gm_n2675, gm_n2676, gm_n2677, gm_n2678, gm_n2679, gm_n268, gm_n2680, gm_n2681, gm_n2682, gm_n2683, gm_n2684, gm_n2685, gm_n2686, gm_n2687, gm_n2688, gm_n2689, gm_n269, gm_n2690, gm_n2691, gm_n2692, gm_n2693, gm_n2694, gm_n2695, gm_n2696, gm_n2697, gm_n2698, gm_n2699, gm_n270, gm_n2700, gm_n2701, gm_n2702, gm_n2703, gm_n2704, gm_n2705, gm_n2706, gm_n2707, gm_n2708, gm_n2709, gm_n271, gm_n2710, gm_n2711, gm_n2712, gm_n2713, gm_n2714, gm_n2715, gm_n2716, gm_n2717, gm_n2718, gm_n2719, gm_n272, gm_n2720, gm_n2721, gm_n2722, gm_n2723, gm_n2724, gm_n2725, gm_n2726, gm_n2727, gm_n2728, gm_n2729, gm_n273, gm_n2730, gm_n2731, gm_n2732, gm_n2733, gm_n2734, gm_n2735, gm_n2736, gm_n2737, gm_n2738, gm_n2739, gm_n274, gm_n2740, gm_n2741, gm_n2742, gm_n2743, gm_n2744, gm_n2745, gm_n2746, gm_n2747, gm_n2748, gm_n275, gm_n2750, gm_n2751, gm_n2752, gm_n2753, gm_n2754, gm_n2755, gm_n2756, gm_n2757, gm_n2758, gm_n2759, gm_n276, gm_n2760, gm_n2761, gm_n2762, gm_n2763, gm_n2764, gm_n2765, gm_n2766, gm_n2767, gm_n2768, gm_n2769, gm_n277, gm_n2770, gm_n2771, gm_n2772, gm_n2773, gm_n2774, gm_n2775, gm_n2776, gm_n2777, gm_n2778, gm_n2779, gm_n278, gm_n2780, gm_n2781, gm_n2782, gm_n2783, gm_n2784, gm_n2785, gm_n2786, gm_n2787, gm_n2788, gm_n2789, gm_n279, gm_n2790, gm_n2791, gm_n2792, gm_n2793, gm_n2794, gm_n2795, gm_n2796, gm_n2797, gm_n2798, gm_n2799, gm_n280, gm_n2800, gm_n2801, gm_n2802, gm_n2803, gm_n2804, gm_n2805, gm_n2806, gm_n2807, gm_n2808, gm_n2809, gm_n281, gm_n2810, gm_n2811, gm_n2812, gm_n2813, gm_n2814, gm_n2815, gm_n2816, gm_n2817, gm_n2818, gm_n2819, gm_n282, gm_n2820, gm_n2821, gm_n2822, gm_n2823, gm_n2824, gm_n2825, gm_n2826, gm_n2827, gm_n2828, gm_n2829, gm_n283, gm_n2830, gm_n2831, gm_n2832, gm_n2833, gm_n2834, gm_n2835, gm_n2836, gm_n2837, gm_n2838, gm_n2839, gm_n284, gm_n2840, gm_n2841, gm_n2842, gm_n2843, gm_n2844, gm_n2845, gm_n2846, gm_n2847, gm_n2848, gm_n2849, gm_n285, gm_n2850, gm_n2851, gm_n2852, gm_n2853, gm_n2854, gm_n2855, gm_n2856, gm_n2857, gm_n2858, gm_n2859, gm_n286, gm_n2860, gm_n2861, gm_n2862, gm_n2863, gm_n2864, gm_n2865, gm_n2866, gm_n2867, gm_n2868, gm_n2869, gm_n287, gm_n2870, gm_n2871, gm_n2872, gm_n2873, gm_n2874, gm_n2875, gm_n2876, gm_n2877, gm_n2878, gm_n2879, gm_n288, gm_n2880, gm_n2881, gm_n2882, gm_n2883, gm_n2884, gm_n2885, gm_n2886, gm_n2887, gm_n2888, gm_n2889, gm_n289, gm_n2890, gm_n2891, gm_n2892, gm_n2893, gm_n2894, gm_n2895, gm_n2896, gm_n2897, gm_n2898, gm_n2899, gm_n290, gm_n2900, gm_n2901, gm_n2902, gm_n2903, gm_n2904, gm_n2905, gm_n2906, gm_n2907, gm_n2908, gm_n2909, gm_n291, gm_n2910, gm_n2911, gm_n2912, gm_n2913, gm_n2914, gm_n2915, gm_n2916, gm_n2917, gm_n2918, gm_n2919, gm_n292, gm_n2920, gm_n2921, gm_n2922, gm_n2923, gm_n2924, gm_n2925, gm_n2926, gm_n2927, gm_n2928, gm_n2929, gm_n293, gm_n2930, gm_n2931, gm_n2932, gm_n2933, gm_n2934, gm_n2935, gm_n2936, gm_n2937, gm_n2938, gm_n2939, gm_n294, gm_n2940, gm_n2941, gm_n2942, gm_n2943, gm_n2944, gm_n2945, gm_n2946, gm_n2947, gm_n2948, gm_n2949, gm_n295, gm_n2950, gm_n2951, gm_n2952, gm_n2953, gm_n2954, gm_n2955, gm_n2956, gm_n2957, gm_n2958, gm_n2959, gm_n296, gm_n2960, gm_n2961, gm_n2962, gm_n2963, gm_n2964, gm_n2965, gm_n2966, gm_n2967, gm_n2968, gm_n2969, gm_n297, gm_n2970, gm_n2971, gm_n2972, gm_n2973, gm_n2974, gm_n2975, gm_n2976, gm_n2977, gm_n2978, gm_n2979, gm_n298, gm_n2980, gm_n2981, gm_n2982, gm_n2983, gm_n2984, gm_n2985, gm_n2986, gm_n2987, gm_n2988, gm_n2989, gm_n299, gm_n2990, gm_n2991, gm_n2992, gm_n2993, gm_n2994, gm_n2995, gm_n2996, gm_n2997, gm_n2998, gm_n2999, gm_n300, gm_n3000, gm_n3001, gm_n3002, gm_n3003, gm_n3004, gm_n3005, gm_n3006, gm_n3007, gm_n3008, gm_n3009, gm_n301, gm_n3010, gm_n3011, gm_n3012, gm_n3013, gm_n3014, gm_n3015, gm_n3016, gm_n3017, gm_n3018, gm_n3019, gm_n302, gm_n3020, gm_n3021, gm_n3022, gm_n3023, gm_n3024, gm_n3025, gm_n3026, gm_n3027, gm_n3028, gm_n3029, gm_n303, gm_n3030, gm_n3031, gm_n3032, gm_n3033, gm_n3034, gm_n3035, gm_n3036, gm_n3037, gm_n3038, gm_n3039, gm_n304, gm_n3040, gm_n3041, gm_n3042, gm_n3043, gm_n3044, gm_n3045, gm_n3046, gm_n3047, gm_n3048, gm_n3049, gm_n305, gm_n3050, gm_n3051, gm_n3052, gm_n3053, gm_n3054, gm_n3055, gm_n3056, gm_n3057, gm_n3058, gm_n3059, gm_n306, gm_n3060, gm_n3061, gm_n3062, gm_n3063, gm_n3064, gm_n3065, gm_n3066, gm_n3067, gm_n3068, gm_n3069, gm_n307, gm_n3070, gm_n3071, gm_n3072, gm_n3073, gm_n3074, gm_n3075, gm_n3076, gm_n3077, gm_n3078, gm_n3079, gm_n308, gm_n3080, gm_n3081, gm_n3082, gm_n3083, gm_n3084, gm_n3085, gm_n3086, gm_n3087, gm_n3088, gm_n3089, gm_n309, gm_n3090, gm_n3091, gm_n3092, gm_n3093, gm_n3094, gm_n3095, gm_n3096, gm_n3097, gm_n3098, gm_n3099, gm_n310, gm_n3100, gm_n3101, gm_n3102, gm_n3103, gm_n3104, gm_n3105, gm_n3106, gm_n3107, gm_n3108, gm_n3109, gm_n311, gm_n3110, gm_n3111, gm_n3112, gm_n3113, gm_n3114, gm_n3115, gm_n3116, gm_n3117, gm_n3118, gm_n3119, gm_n312, gm_n3120, gm_n3121, gm_n3122, gm_n3123, gm_n3124, gm_n3125, gm_n3126, gm_n3127, gm_n3128, gm_n3129, gm_n313, gm_n3130, gm_n3131, gm_n3132, gm_n3133, gm_n3134, gm_n3135, gm_n3136, gm_n3137, gm_n3138, gm_n3139, gm_n314, gm_n3140, gm_n3141, gm_n3142, gm_n3143, gm_n3144, gm_n3145, gm_n3146, gm_n3147, gm_n3148, gm_n3149, gm_n315, gm_n3150, gm_n3151, gm_n3152, gm_n3153, gm_n3154, gm_n3155, gm_n3156, gm_n3157, gm_n3158, gm_n3159, gm_n316, gm_n3160, gm_n3161, gm_n3162, gm_n3163, gm_n3164, gm_n3165, gm_n3166, gm_n3167, gm_n3168, gm_n3169, gm_n317, gm_n3170, gm_n3171, gm_n3172, gm_n3173, gm_n3174, gm_n3175, gm_n3176, gm_n3177, gm_n3178, gm_n3179, gm_n318, gm_n3180, gm_n3181, gm_n3182, gm_n3183, gm_n3184, gm_n3185, gm_n3186, gm_n3187, gm_n3188, gm_n3189, gm_n319, gm_n3190, gm_n3191, gm_n3192, gm_n3193, gm_n3194, gm_n3195, gm_n3196, gm_n3197, gm_n3198, gm_n3199, gm_n320, gm_n3200, gm_n3201, gm_n3202, gm_n3203, gm_n3204, gm_n3205, gm_n3206, gm_n3207, gm_n3208, gm_n3209, gm_n321, gm_n3210, gm_n3211, gm_n3212, gm_n3213, gm_n3214, gm_n3215, gm_n3216, gm_n3217, gm_n3218, gm_n3219, gm_n322, gm_n3220, gm_n3221, gm_n3222, gm_n3223, gm_n3224, gm_n3225, gm_n3226, gm_n3227, gm_n3228, gm_n3229, gm_n323, gm_n3230, gm_n3231, gm_n3232, gm_n3233, gm_n3234, gm_n3235, gm_n3236, gm_n3237, gm_n3238, gm_n3239, gm_n324, gm_n3240, gm_n3241, gm_n3242, gm_n3243, gm_n3244, gm_n3245, gm_n3246, gm_n3247, gm_n3248, gm_n3249, gm_n325, gm_n3250, gm_n3251, gm_n3252, gm_n3253, gm_n3254, gm_n3255, gm_n3256, gm_n3257, gm_n3258, gm_n3259, gm_n326, gm_n3260, gm_n3261, gm_n3262, gm_n3263, gm_n3264, gm_n3265, gm_n3266, gm_n3267, gm_n3268, gm_n3269, gm_n327, gm_n3270, gm_n3271, gm_n3272, gm_n3273, gm_n3274, gm_n3275, gm_n3276, gm_n3277, gm_n3278, gm_n3279, gm_n328, gm_n3280, gm_n3281, gm_n3282, gm_n3283, gm_n3284, gm_n3285, gm_n3286, gm_n3287, gm_n3288, gm_n3289, gm_n329, gm_n3290, gm_n3291, gm_n3292, gm_n3293, gm_n3294, gm_n3295, gm_n3296, gm_n3297, gm_n3298, gm_n3299, gm_n330, gm_n3300, gm_n3301, gm_n3302, gm_n3303, gm_n3304, gm_n3305, gm_n3306, gm_n3307, gm_n3308, gm_n3309, gm_n331, gm_n3310, gm_n3311, gm_n3312, gm_n3313, gm_n3314, gm_n3315, gm_n3316, gm_n3317, gm_n3318, gm_n3319, gm_n332, gm_n3320, gm_n3321, gm_n3322, gm_n3323, gm_n3324, gm_n3325, gm_n3326, gm_n3327, gm_n3328, gm_n3329, gm_n333, gm_n3330, gm_n3331, gm_n3332, gm_n3333, gm_n3334, gm_n3335, gm_n3336, gm_n3337, gm_n3338, gm_n3339, gm_n334, gm_n3340, gm_n3341, gm_n3342, gm_n3343, gm_n3344, gm_n3345, gm_n3346, gm_n3347, gm_n3348, gm_n3349, gm_n335, gm_n3350, gm_n3351, gm_n3352, gm_n3353, gm_n3354, gm_n3355, gm_n3356, gm_n3357, gm_n3358, gm_n3359, gm_n336, gm_n3360, gm_n3361, gm_n3362, gm_n3363, gm_n3364, gm_n3365, gm_n3366, gm_n3367, gm_n3368, gm_n3369, gm_n337, gm_n3370, gm_n3371, gm_n3372, gm_n3373, gm_n3374, gm_n3375, gm_n3376, gm_n3377, gm_n3378, gm_n3379, gm_n338, gm_n3380, gm_n3381, gm_n3382, gm_n3383, gm_n3384, gm_n3385, gm_n3386, gm_n3387, gm_n3388, gm_n3389, gm_n339, gm_n3390, gm_n3391, gm_n3392, gm_n3393, gm_n3394, gm_n3395, gm_n3396, gm_n3397, gm_n3398, gm_n3399, gm_n340, gm_n3400, gm_n3401, gm_n3402, gm_n3403, gm_n3404, gm_n3405, gm_n3406, gm_n3407, gm_n3408, gm_n3409, gm_n341, gm_n3410, gm_n3411, gm_n3412, gm_n3413, gm_n3414, gm_n3415, gm_n3416, gm_n3417, gm_n3418, gm_n3419, gm_n342, gm_n3420, gm_n3421, gm_n3422, gm_n3423, gm_n3424, gm_n3425, gm_n3426, gm_n3427, gm_n3428, gm_n3429, gm_n343, gm_n3430, gm_n3431, gm_n3432, gm_n3433, gm_n3434, gm_n3435, gm_n3436, gm_n3437, gm_n3438, gm_n3439, gm_n344, gm_n3440, gm_n3441, gm_n3442, gm_n3443, gm_n3444, gm_n3445, gm_n3446, gm_n3447, gm_n3448, gm_n3449, gm_n345, gm_n3450, gm_n3451, gm_n3452, gm_n3453, gm_n3454, gm_n3455, gm_n3456, gm_n3457, gm_n3458, gm_n3459, gm_n346, gm_n3460, gm_n3461, gm_n3462, gm_n3463, gm_n3464, gm_n3465, gm_n3466, gm_n347, gm_n348, gm_n349, gm_n350, gm_n351, gm_n352, gm_n353, gm_n354, gm_n355, gm_n356, gm_n357, gm_n358, gm_n359, gm_n360, gm_n361, gm_n362, gm_n363, gm_n364, gm_n365, gm_n366, gm_n367, gm_n368, gm_n369, gm_n370, gm_n371, gm_n372, gm_n373, gm_n374, gm_n375, gm_n376, gm_n377, gm_n378, gm_n379, gm_n380, gm_n381, gm_n382, gm_n383, gm_n384, gm_n385, gm_n386, gm_n387, gm_n388, gm_n389, gm_n390, gm_n391, gm_n392, gm_n393, gm_n394, gm_n395, gm_n396, gm_n397, gm_n398, gm_n399, gm_n400, gm_n401, gm_n402, gm_n403, gm_n404, gm_n405, gm_n406, gm_n407, gm_n408, gm_n409, gm_n410, gm_n411, gm_n412, gm_n413, gm_n414, gm_n415, gm_n416, gm_n417, gm_n418, gm_n419, gm_n420, gm_n421, gm_n422, gm_n423, gm_n424, gm_n425, gm_n426, gm_n427, gm_n428, gm_n429, gm_n430, gm_n431, gm_n432, gm_n433, gm_n434, gm_n435, gm_n436, gm_n437, gm_n438, gm_n439, gm_n440, gm_n441, gm_n442, gm_n443, gm_n444, gm_n445, gm_n446, gm_n447, gm_n448, gm_n449, gm_n450, gm_n451, gm_n452, gm_n453, gm_n454, gm_n455, gm_n456, gm_n457, gm_n458, gm_n459, gm_n460, gm_n461, gm_n462, gm_n463, gm_n464, gm_n465, gm_n466, gm_n467, gm_n468, gm_n469, gm_n470, gm_n471, gm_n472, gm_n473, gm_n474, gm_n475, gm_n476, gm_n477, gm_n478, gm_n479, gm_n480, gm_n481, gm_n482, gm_n483, gm_n484, gm_n485, gm_n486, gm_n487, gm_n488, gm_n489, gm_n490, gm_n491, gm_n492, gm_n493, gm_n494, gm_n495, gm_n496, gm_n497, gm_n498, gm_n499, gm_n500, gm_n501, gm_n502, gm_n503, gm_n504, gm_n505, gm_n506, gm_n508, gm_n509, gm_n510, gm_n511, gm_n512, gm_n513, gm_n514, gm_n515, gm_n516, gm_n517, gm_n518, gm_n519, gm_n520, gm_n521, gm_n522, gm_n523, gm_n524, gm_n525, gm_n526, gm_n527, gm_n528, gm_n529, gm_n530, gm_n531, gm_n532, gm_n533, gm_n534, gm_n535, gm_n536, gm_n537, gm_n538, gm_n539, gm_n54, gm_n540, gm_n541, gm_n542, gm_n543, gm_n544, gm_n545, gm_n546, gm_n547, gm_n548, gm_n549, gm_n55, gm_n550, gm_n551, gm_n552, gm_n553, gm_n554, gm_n555, gm_n556, gm_n557, gm_n558, gm_n559, gm_n56, gm_n560, gm_n561, gm_n562, gm_n563, gm_n564, gm_n565, gm_n566, gm_n567, gm_n568, gm_n569, gm_n57, gm_n570, gm_n571, gm_n572, gm_n573, gm_n574, gm_n575, gm_n576, gm_n577, gm_n578, gm_n579, gm_n58, gm_n580, gm_n581, gm_n582, gm_n583, gm_n584, gm_n585, gm_n586, gm_n587, gm_n588, gm_n589, gm_n59, gm_n590, gm_n591, gm_n592, gm_n593, gm_n594, gm_n595, gm_n596, gm_n597, gm_n598, gm_n599, gm_n60, gm_n600, gm_n601, gm_n602, gm_n603, gm_n604, gm_n605, gm_n606, gm_n607, gm_n608, gm_n609, gm_n61, gm_n610, gm_n611, gm_n612, gm_n613, gm_n614, gm_n615, gm_n616, gm_n617, gm_n618, gm_n619, gm_n62, gm_n620, gm_n621, gm_n622, gm_n623, gm_n624, gm_n625, gm_n626, gm_n627, gm_n628, gm_n629, gm_n63, gm_n630, gm_n631, gm_n632, gm_n633, gm_n634, gm_n635, gm_n636, gm_n637, gm_n638, gm_n639, gm_n64, gm_n640, gm_n641, gm_n642, gm_n643, gm_n644, gm_n645, gm_n646, gm_n647, gm_n648, gm_n649, gm_n65, gm_n650, gm_n651, gm_n652, gm_n653, gm_n654, gm_n655, gm_n656, gm_n657, gm_n658, gm_n659, gm_n66, gm_n660, gm_n661, gm_n662, gm_n663, gm_n664, gm_n665, gm_n666, gm_n667, gm_n668, gm_n669, gm_n67, gm_n670, gm_n671, gm_n672, gm_n673, gm_n674, gm_n675, gm_n676, gm_n677, gm_n678, gm_n679, gm_n68, gm_n680, gm_n681, gm_n682, gm_n683, gm_n684, gm_n685, gm_n686, gm_n687, gm_n688, gm_n689, gm_n69, gm_n690, gm_n691, gm_n692, gm_n693, gm_n694, gm_n695, gm_n696, gm_n697, gm_n698, gm_n699, gm_n70, gm_n700, gm_n701, gm_n702, gm_n703, gm_n704, gm_n705, gm_n706, gm_n707, gm_n708, gm_n709, gm_n71, gm_n710, gm_n711, gm_n712, gm_n713, gm_n714, gm_n715, gm_n716, gm_n717, gm_n718, gm_n719, gm_n72, gm_n720, gm_n721, gm_n722, gm_n723, gm_n724, gm_n725, gm_n726, gm_n727, gm_n728, gm_n729, gm_n73, gm_n730, gm_n731, gm_n732, gm_n733, gm_n734, gm_n735, gm_n736, gm_n737, gm_n738, gm_n739, gm_n74, gm_n740, gm_n741, gm_n742, gm_n743, gm_n744, gm_n745, gm_n746, gm_n747, gm_n748, gm_n749, gm_n75, gm_n750, gm_n751, gm_n752, gm_n753, gm_n754, gm_n755, gm_n756, gm_n757, gm_n758, gm_n759, gm_n76, gm_n760, gm_n761, gm_n762, gm_n763, gm_n764, gm_n765, gm_n766, gm_n767, gm_n768, gm_n769, gm_n77, gm_n770, gm_n771, gm_n772, gm_n774, gm_n775, gm_n776, gm_n777, gm_n778, gm_n779, gm_n78, gm_n780, gm_n781, gm_n782, gm_n783, gm_n784, gm_n785, gm_n786, gm_n787, gm_n788, gm_n789, gm_n79, gm_n790, gm_n791, gm_n792, gm_n793, gm_n794, gm_n795, gm_n796, gm_n797, gm_n798, gm_n799, gm_n80, gm_n800, gm_n801, gm_n802, gm_n803, gm_n804, gm_n805, gm_n806, gm_n807, gm_n808, gm_n809, gm_n81, gm_n810, gm_n811, gm_n812, gm_n813, gm_n814, gm_n815, gm_n816, gm_n817, gm_n818, gm_n819, gm_n82, gm_n820, gm_n821, gm_n822, gm_n823, gm_n824, gm_n825, gm_n826, gm_n827, gm_n828, gm_n829, gm_n83, gm_n830, gm_n831, gm_n832, gm_n833, gm_n834, gm_n835, gm_n836, gm_n837, gm_n838, gm_n839, gm_n84, gm_n840, gm_n841, gm_n842, gm_n843, gm_n844, gm_n845, gm_n846, gm_n847, gm_n848, gm_n849, gm_n85, gm_n850, gm_n851, gm_n852, gm_n853, gm_n854, gm_n855, gm_n856, gm_n857, gm_n858, gm_n859, gm_n86, gm_n860, gm_n861, gm_n862, gm_n863, gm_n864, gm_n865, gm_n866, gm_n867, gm_n868, gm_n869, gm_n87, gm_n870, gm_n871, gm_n872, gm_n873, gm_n874, gm_n875, gm_n876, gm_n877, gm_n878, gm_n879, gm_n88, gm_n880, gm_n881, gm_n882, gm_n883, gm_n884, gm_n885, gm_n886, gm_n887, gm_n888, gm_n889, gm_n89, gm_n890, gm_n891, gm_n892, gm_n893, gm_n894, gm_n895, gm_n896, gm_n897, gm_n898, gm_n899, gm_n90, gm_n900, gm_n901, gm_n902, gm_n903, gm_n904, gm_n905, gm_n906, gm_n907, gm_n908, gm_n909, gm_n91, gm_n910, gm_n911, gm_n912, gm_n913, gm_n914, gm_n915, gm_n916, gm_n917, gm_n918, gm_n919, gm_n92, gm_n920, gm_n921, gm_n922, gm_n923, gm_n924, gm_n925, gm_n926, gm_n927, gm_n928, gm_n929, gm_n93, gm_n930, gm_n931, gm_n932, gm_n933, gm_n934, gm_n935, gm_n936, gm_n937, gm_n938, gm_n939, gm_n94, gm_n940, gm_n941, gm_n942, gm_n943, gm_n944, gm_n945, gm_n946, gm_n947, gm_n948, gm_n949, gm_n95, gm_n950, gm_n951, gm_n952, gm_n953, gm_n954, gm_n955, gm_n956, gm_n957, gm_n958, gm_n959, gm_n96, gm_n960, gm_n961, gm_n962, gm_n963, gm_n964, gm_n965, gm_n966, gm_n967, gm_n968, gm_n969, gm_n97, gm_n970, gm_n971, gm_n972, gm_n973, gm_n974, gm_n975, gm_n976, gm_n977, gm_n978, gm_n979, gm_n98, gm_n980, gm_n981, gm_n982, gm_n983, gm_n984, gm_n985, gm_n986, gm_n987, gm_n988, gm_n989, gm_n99, gm_n991, gm_n992, gm_n993, gm_n994, gm_n995, gm_n996, gm_n997, gm_n998, gm_n999;
	wire t_3, t_1, t_0, t_2;
	not (gm_n54, in_27);
	not (gm_n55, in_31);
	and (gm_n56, in_30, in_29, in_28);
	not (gm_n57, gm_n56);
	not (gm_n58, in_19);
	not (gm_n59, in_26);
	nor (gm_n60, gm_n59, in_25, in_24);
	not (gm_n61, in_11);
	not (gm_n62, in_15);
	not (gm_n63, in_12);
	not (gm_n64, in_14);
	nor (gm_n65, gm_n64, in_13, gm_n63);
	not (gm_n66, in_10);
	not (gm_n67, in_1);
	not (gm_n68, in_3);
	nor (gm_n69, in_2, gm_n67, in_0, in_4, gm_n68);
	not (gm_n70, in_5);
	nor (gm_n71, in_7, in_6, gm_n70);
	and (gm_n72, gm_n66, in_9, in_8, gm_n71, gm_n69);
	not (gm_n73, in_16);
	nor (gm_n74, in_18, in_17, gm_n73);
	and (gm_n75, gm_n65, gm_n62, gm_n61, gm_n74, gm_n72);
	not (gm_n76, in_20);
	nor (gm_n77, in_22, in_21, gm_n76);
	nand (gm_n78, gm_n60, in_23, gm_n58, gm_n77, gm_n75);
	nor (gm_n79, gm_n57, gm_n55, gm_n54, gm_n78);
	not (gm_n80, in_29);
	nor (gm_n81, gm_n55, in_30, gm_n80);
	not (gm_n82, in_24);
	not (gm_n83, in_28);
	nor (gm_n84, in_27, in_26, in_25);
	not (gm_n85, gm_n84);
	not (gm_n86, in_21);
	not (gm_n87, in_22);
	nor (gm_n88, in_23, gm_n87, gm_n86);
	not (gm_n89, gm_n88);
	nor (gm_n90, in_19, in_18, in_17);
	and (gm_n91, in_15, in_14, in_13);
	nand (gm_n92, gm_n61, gm_n66, in_9);
	nand (gm_n93, in_7, in_6, gm_n70);
	not (gm_n94, in_0);
	nand (gm_n95, in_2, gm_n67, gm_n94, in_4, in_3);
	nor (gm_n96, gm_n92, in_12, in_8, gm_n95, gm_n93);
	nand (gm_n97, gm_n90, gm_n76, gm_n73, gm_n96, gm_n91);
	nor (gm_n98, gm_n85, gm_n83, gm_n82, gm_n97, gm_n89);
	nand (gm_n99, gm_n98, gm_n81);
	not (gm_n100, in_30);
	nor (gm_n101, gm_n55, gm_n100, in_29);
	nor (gm_n102, in_27, gm_n59, in_25);
	and (gm_n103, in_23, in_22, in_21);
	not (gm_n104, gm_n103);
	not (gm_n105, in_17);
	not (gm_n106, in_18);
	nor (gm_n107, in_19, gm_n106, gm_n105);
	not (gm_n108, gm_n107);
	nand (gm_n109, gm_n62, gm_n64, in_13);
	nor (gm_n110, gm_n61, gm_n66, in_9);
	not (gm_n111, gm_n110);
	not (gm_n112, in_2);
	not (gm_n113, in_4);
	nand (gm_n114, gm_n112, gm_n67, gm_n94, gm_n113, in_3);
	not (gm_n115, in_6);
	nand (gm_n116, in_7, gm_n115, in_5);
	or (gm_n117, gm_n116, gm_n114);
	or (gm_n118, gm_n109, in_12, in_8, gm_n117, gm_n111);
	nor (gm_n119, gm_n104, in_20, gm_n73, gm_n118, gm_n108);
	nand (gm_n120, gm_n101, gm_n83, in_24, gm_n119, gm_n102);
	nor (gm_n121, gm_n106, in_17, in_16);
	not (gm_n122, gm_n121);
	nor (gm_n123, gm_n64, in_13, in_12);
	not (gm_n124, in_8);
	nand (gm_n125, in_10, in_9, gm_n124);
	not (gm_n126, gm_n125);
	nor (gm_n127, in_7, gm_n115, in_5);
	nor (gm_n128, in_2, gm_n67, gm_n94, gm_n113, gm_n68);
	nand (gm_n129, gm_n126, gm_n123, in_11, gm_n128, gm_n127);
	nor (gm_n130, in_22, gm_n86, in_20);
	not (gm_n131, gm_n130);
	nor (gm_n132, gm_n122, in_19, gm_n62, gm_n131, gm_n129);
	not (gm_n133, in_25);
	nor (gm_n134, in_26, gm_n133, gm_n82);
	nand (gm_n135, gm_n56, in_27, in_23, gm_n134, gm_n132);
	nor (gm_n136, gm_n135, gm_n55);
	nor (gm_n137, in_31, in_30, in_29);
	not (gm_n138, gm_n137);
	nor (gm_n139, gm_n54, in_26, in_25);
	not (gm_n140, gm_n139);
	nor (gm_n141, gm_n58, gm_n106, in_17);
	nor (gm_n142, in_15, in_14, in_13);
	not (gm_n143, gm_n142);
	and (gm_n144, in_7, in_6, in_5);
	and (gm_n145, in_2, in_1, in_0);
	nand (gm_n146, gm_n144, gm_n113, gm_n68, gm_n145);
	nor (gm_n147, gm_n92, in_12, in_8, gm_n146, gm_n143);
	nand (gm_n148, gm_n103, in_20, in_16, gm_n147, gm_n141);
	nor (gm_n149, gm_n138, in_28, in_24, gm_n148, gm_n140);
	nor (gm_n150, gm_n62, gm_n64, in_13);
	not (gm_n151, in_7);
	nand (gm_n152, gm_n151, gm_n115, in_5);
	and (gm_n153, in_11, in_10, in_9);
	not (gm_n154, gm_n153);
	nor (gm_n155, gm_n152, gm_n63, in_8, gm_n154, gm_n95);
	nand (gm_n156, gm_n150, in_17, in_16, gm_n155);
	nand (gm_n157, in_20, in_19, gm_n106);
	not (gm_n158, in_23);
	nor (gm_n159, gm_n82, gm_n158, in_22);
	not (gm_n160, gm_n159);
	nor (gm_n161, gm_n156, gm_n133, gm_n86, gm_n160, gm_n157);
	nor (gm_n162, in_28, in_27, gm_n59);
	nand (gm_n163, gm_n55, gm_n100, gm_n80, gm_n162, gm_n161);
	nor (gm_n164, gm_n58, in_18, in_17);
	not (gm_n165, gm_n164);
	nor (gm_n166, gm_n62, in_14, in_13);
	nor (gm_n167, in_11, in_10, in_9);
	nand (gm_n168, in_2, in_1, gm_n94, in_4, in_3);
	nor (gm_n169, gm_n168, gm_n93, in_8);
	nand (gm_n170, gm_n166, gm_n73, in_12, gm_n169, gm_n167);
	nor (gm_n171, gm_n89, in_24, gm_n76, gm_n170, gm_n165);
	nand (gm_n172, gm_n102, gm_n81, in_28, gm_n171);
	nor (gm_n173, in_22, gm_n86, gm_n76);
	nor (gm_n174, gm_n106, in_17, gm_n73);
	not (gm_n175, in_13);
	nor (gm_n176, gm_n62, in_14, gm_n175);
	not (gm_n177, gm_n176);
	nand (gm_n178, in_2, in_1, gm_n94, gm_n113, gm_n68);
	or (gm_n179, gm_n152, in_12, in_8, gm_n178, gm_n154);
	nor (gm_n180, gm_n179, gm_n177);
	nand (gm_n181, gm_n173, in_23, in_19, gm_n180, gm_n174);
	nor (gm_n182, gm_n59, gm_n133, in_24);
	not (gm_n183, gm_n182);
	nor (gm_n184, gm_n57, in_31, gm_n54, gm_n183, gm_n181);
	not (gm_n185, gm_n101);
	nor (gm_n186, in_27, gm_n59, gm_n133);
	not (gm_n187, gm_n141);
	nand (gm_n188, gm_n62, in_14, in_13);
	nor (gm_n189, gm_n151, in_6, gm_n70);
	nand (gm_n190, gm_n69, in_12, in_8, gm_n189, gm_n110);
	nor (gm_n191, gm_n187, in_20, gm_n73, gm_n190, gm_n188);
	nor (gm_n192, in_23, in_22, gm_n86);
	nand (gm_n193, gm_n186, gm_n83, gm_n82, gm_n192, gm_n191);
	nor (gm_n194, gm_n193, gm_n185);
	nand (gm_n195, gm_n55, gm_n100, in_29);
	not (gm_n196, gm_n195);
	not (gm_n197, gm_n90);
	not (gm_n198, in_9);
	nor (gm_n199, in_11, in_10, gm_n198);
	nor (gm_n200, in_15, in_14, gm_n175);
	and (gm_n201, gm_n127, gm_n69, gm_n124);
	nand (gm_n202, gm_n199, in_16, gm_n63, gm_n201, gm_n200);
	nor (gm_n203, gm_n89, in_24, gm_n76, gm_n202, gm_n197);
	nand (gm_n204, gm_n196, gm_n84, gm_n83, gm_n203);
	nor (gm_n205, gm_n158, gm_n87, in_21);
	not (gm_n206, gm_n205);
	nor (gm_n207, in_15, gm_n64, in_13);
	nor (gm_n208, gm_n112, in_1, gm_n94, gm_n113, in_3);
	and (gm_n209, gm_n144, in_12, in_8, gm_n208, gm_n153);
	nand (gm_n210, gm_n141, gm_n76, gm_n73, gm_n209, gm_n207);
	nor (gm_n211, gm_n140, in_28, gm_n82, gm_n210, gm_n206);
	nand (gm_n212, gm_n211, gm_n137);
	nor (gm_n213, in_31, gm_n100, in_29);
	not (gm_n214, gm_n213);
	and (gm_n215, in_27, in_26, in_25);
	not (gm_n216, gm_n215);
	nor (gm_n217, gm_n158, in_22, gm_n86);
	nor (gm_n218, gm_n151, gm_n115, in_5);
	nor (gm_n219, gm_n112, in_1, in_0, in_4, gm_n68);
	and (gm_n220, gm_n219, gm_n218, gm_n124);
	and (gm_n221, gm_n110, in_16, in_12, gm_n220, gm_n142);
	nand (gm_n222, gm_n90, in_24, gm_n76, gm_n221, gm_n217);
	nor (gm_n223, gm_n216, gm_n214, gm_n83, gm_n222);
	not (gm_n224, gm_n102);
	nor (gm_n225, gm_n55, in_30, in_29);
	not (gm_n226, gm_n225);
	nor (gm_n227, gm_n158, in_22, in_21);
	nor (gm_n228, in_11, gm_n66, gm_n198);
	nand (gm_n229, in_2, gm_n67, gm_n94, in_4, gm_n68);
	nor (gm_n230, gm_n151, gm_n115, gm_n70, gm_n229, gm_n124);
	and (gm_n231, gm_n207, in_16, in_12, gm_n230, gm_n228);
	nand (gm_n232, gm_n164, in_24, in_20, gm_n231, gm_n227);
	nor (gm_n233, gm_n226, gm_n224, gm_n83, gm_n232);
	not (gm_n234, gm_n81);
	nor (gm_n235, in_19, gm_n106, in_17);
	not (gm_n236, gm_n166);
	nand (gm_n237, gm_n61, in_10, gm_n198);
	nand (gm_n238, in_8, gm_n113, gm_n68, gm_n145, gm_n127);
	nor (gm_n239, gm_n236, gm_n73, gm_n63, gm_n238, gm_n237);
	nand (gm_n240, gm_n217, in_24, gm_n76, gm_n239, gm_n235);
	nor (gm_n241, gm_n85, gm_n234, in_28, gm_n240);
	nor (gm_n242, in_11, gm_n66, in_9);
	nor (gm_n243, in_2, gm_n67, gm_n94, in_4, in_3);
	and (gm_n244, gm_n144, gm_n63, gm_n124, gm_n243, gm_n242);
	and (gm_n245, gm_n107, gm_n76, in_16, gm_n244, gm_n142);
	nand (gm_n246, gm_n103, in_28, gm_n82, gm_n245, gm_n215);
	nor (gm_n247, gm_n246, gm_n185);
	not (gm_n248, gm_n186);
	not (gm_n249, gm_n91);
	or (gm_n250, gm_n168, gm_n116, gm_n124);
	nor (gm_n251, gm_n249, gm_n73, in_12, gm_n250, gm_n237);
	nand (gm_n252, gm_n107, in_24, gm_n76, gm_n251, gm_n205);
	nor (gm_n253, gm_n248, gm_n185, gm_n83, gm_n252);
	nor (gm_n254, gm_n241, gm_n233, gm_n223, gm_n253, gm_n247);
	nor (gm_n255, in_23, gm_n87, in_21);
	nor (gm_n256, gm_n61, in_10, gm_n198);
	nor (gm_n257, in_2, gm_n67, in_0, in_4, in_3);
	nand (gm_n258, gm_n144, in_12, gm_n124, gm_n257, gm_n256);
	nor (gm_n259, gm_n197, gm_n76, gm_n73, gm_n258, gm_n249);
	nand (gm_n260, gm_n139, in_28, in_24, gm_n259, gm_n255);
	nor (gm_n261, gm_n260, gm_n234);
	nand (gm_n262, gm_n54, gm_n59, in_25);
	nor (gm_n263, in_23, in_22, in_21);
	nor (gm_n264, gm_n151, in_6, in_5);
	nor (gm_n265, in_2, gm_n67, in_0, gm_n113, in_3);
	nand (gm_n266, gm_n265, gm_n264, gm_n124);
	nor (gm_n267, gm_n177, gm_n73, in_12, gm_n266, gm_n237);
	nand (gm_n268, gm_n235, gm_n82, gm_n76, gm_n267, gm_n263);
	nor (gm_n269, gm_n262, gm_n234, gm_n83, gm_n268);
	nor (gm_n270, gm_n58, in_18, gm_n105);
	nand (gm_n271, in_2, in_1, gm_n94, in_4, gm_n68);
	nor (gm_n272, gm_n271, gm_n152, in_8);
	and (gm_n273, gm_n200, in_16, gm_n63, gm_n272, gm_n167);
	nand (gm_n274, gm_n103, in_24, gm_n76, gm_n273, gm_n270);
	nor (gm_n275, gm_n195, gm_n248, gm_n83, gm_n274);
	nor (gm_n276, gm_n275, gm_n269, gm_n261);
	nand (gm_n277, gm_n112, in_1, gm_n94, gm_n113, gm_n68);
	nor (gm_n278, gm_n277, gm_n152, gm_n124);
	and (gm_n279, gm_n166, in_16, gm_n63, gm_n278, gm_n242);
	nand (gm_n280, gm_n141, in_24, in_20, gm_n279, gm_n227);
	nor (gm_n281, gm_n216, gm_n185, in_28, gm_n280);
	nand (gm_n282, in_11, gm_n66, in_9);
	nor (gm_n283, in_2, in_1, in_0, gm_n113, gm_n68);
	nand (gm_n284, gm_n283, gm_n144);
	nor (gm_n285, gm_n177, in_12, gm_n124, gm_n284, gm_n282);
	nand (gm_n286, gm_n205, gm_n76, in_16, gm_n285, gm_n235);
	nor (gm_n287, gm_n140, in_28, gm_n82, gm_n286, gm_n214);
	nand (gm_n288, in_11, gm_n66, gm_n198);
	and (gm_n289, gm_n145, in_4, gm_n68);
	nand (gm_n290, gm_n289, gm_n218, in_8);
	nor (gm_n291, gm_n188, gm_n73, in_12, gm_n290, gm_n288);
	nand (gm_n292, gm_n217, gm_n82, gm_n76, gm_n291, gm_n270);
	nor (gm_n293, gm_n262, gm_n214, in_28, gm_n292);
	nor (gm_n294, gm_n293, gm_n287, gm_n281);
	nand (gm_n295, gm_n254, gm_n212, gm_n204, gm_n294, gm_n276);
	and (gm_n296, in_22, in_21, in_20);
	not (gm_n297, gm_n296);
	nand (gm_n298, gm_n112, gm_n67, in_0, gm_n113, gm_n68);
	nor (gm_n299, gm_n298, gm_n116);
	nor (gm_n300, gm_n66, in_9, in_8);
	nand (gm_n301, gm_n123, gm_n62, gm_n61, gm_n300, gm_n299);
	nor (gm_n302, in_18, gm_n105, in_16);
	not (gm_n303, gm_n302);
	nor (gm_n304, gm_n297, in_23, gm_n58, gm_n303, gm_n301);
	nor (gm_n305, in_26, in_25, in_24);
	nor (gm_n306, in_30, in_29, in_28);
	nand (gm_n307, gm_n304, in_31, in_27, gm_n306, gm_n305);
	nor (gm_n308, gm_n100, in_29, in_28);
	nor (gm_n309, gm_n59, in_25, gm_n82);
	nor (gm_n310, in_7, in_6, in_5);
	nor (gm_n311, gm_n112, in_1, gm_n94, gm_n113, gm_n68);
	nand (gm_n312, gm_n311, gm_n310);
	and (gm_n313, in_14, in_13, in_12);
	not (gm_n314, gm_n313);
	or (gm_n315, gm_n125, in_15, in_11, gm_n314, gm_n312);
	nor (gm_n316, gm_n87, gm_n86, in_20);
	not (gm_n317, gm_n316);
	nor (gm_n318, gm_n122, gm_n158, gm_n58, gm_n317, gm_n315);
	nand (gm_n319, gm_n308, gm_n55, in_27, gm_n318, gm_n309);
	nor (gm_n320, in_2, in_1, in_0, in_3);
	nand (gm_n321, gm_n115, in_5, in_4, gm_n320, gm_n151);
	nand (gm_n322, gm_n66, gm_n198, in_8);
	or (gm_n323, gm_n175, in_12, in_11, gm_n322, gm_n321);
	nor (gm_n324, in_16, gm_n62, gm_n64, gm_n323, gm_n105);
	and (gm_n325, in_20, in_19, in_18);
	and (gm_n326, in_24, in_23, in_22);
	and (gm_n327, gm_n324, gm_n133, in_21, gm_n326, gm_n325);
	nor (gm_n328, in_28, in_27, in_26);
	nand (gm_n329, gm_n55, in_30, gm_n80, gm_n328, gm_n327);
	nand (gm_n330, gm_n329, gm_n319, gm_n307);
	not (gm_n331, gm_n174);
	and (gm_n332, gm_n115, gm_n70, in_4, gm_n320, in_7);
	nand (gm_n333, gm_n65, in_15, in_11, gm_n332, gm_n126);
	nor (gm_n334, gm_n87, in_21, gm_n76);
	not (gm_n335, gm_n334);
	nor (gm_n336, gm_n331, gm_n158, in_19, gm_n335, gm_n333);
	nor (gm_n337, gm_n100, gm_n80, in_28);
	nand (gm_n338, gm_n309, in_31, in_27, gm_n337, gm_n336);
	not (gm_n339, gm_n262);
	nor (gm_n340, gm_n61, in_10, in_9);
	and (gm_n341, gm_n219, gm_n71, gm_n124);
	nand (gm_n342, gm_n142, gm_n73, gm_n63, gm_n341, gm_n340);
	nor (gm_n343, gm_n108, gm_n82, in_20, gm_n342, gm_n206);
	nand (gm_n344, gm_n339, gm_n81, gm_n83, gm_n343);
	nand (gm_n345, gm_n151, in_6, in_5);
	nor (gm_n346, gm_n345, gm_n298, in_8);
	nand (gm_n347, gm_n150, in_16, gm_n63, gm_n346, gm_n256);
	nor (gm_n348, gm_n108, gm_n82, gm_n76, gm_n347, gm_n206);
	nand (gm_n349, gm_n139, gm_n137, gm_n83, gm_n348);
	nand (gm_n350, gm_n349, gm_n344, gm_n338);
	nor (gm_n351, gm_n295, gm_n194, gm_n184, gm_n350, gm_n330);
	nand (gm_n352, gm_n61, in_10, in_9);
	nand (gm_n353, gm_n283, gm_n189, in_8);
	nor (gm_n354, gm_n143, in_16, gm_n63, gm_n353, gm_n352);
	nand (gm_n355, gm_n235, in_24, in_20, gm_n354, gm_n263);
	nor (gm_n356, gm_n248, gm_n234, gm_n83, gm_n355);
	not (gm_n357, gm_n308);
	nor (gm_n358, in_22, in_21, in_20);
	nor (gm_n359, in_18, in_17, in_16);
	not (gm_n360, gm_n359);
	nor (gm_n361, in_2, in_1, in_0, in_4, in_3);
	nand (gm_n362, gm_n66, in_9, gm_n124, gm_n361, gm_n310);
	nand (gm_n363, gm_n64, in_13, in_12);
	nor (gm_n364, gm_n360, gm_n62, in_11, gm_n363, gm_n362);
	nand (gm_n365, gm_n60, in_23, gm_n58, gm_n364, gm_n358);
	nor (gm_n366, gm_n357, gm_n55, gm_n54, gm_n365);
	nor (gm_n367, gm_n54, gm_n59, in_25);
	not (gm_n368, gm_n367);
	nand (gm_n369, gm_n128, gm_n71);
	nor (gm_n370, gm_n177, gm_n63, in_8, gm_n369, gm_n352);
	nand (gm_n371, gm_n107, gm_n76, gm_n73, gm_n370, gm_n255);
	nor (gm_n372, gm_n234, in_28, gm_n82, gm_n371, gm_n368);
	nor (gm_n373, gm_n372, gm_n366, gm_n356);
	nand (gm_n374, gm_n62, in_14, gm_n175);
	or (gm_n375, gm_n271, gm_n116, in_8);
	nor (gm_n376, gm_n374, gm_n73, gm_n63, gm_n375, gm_n282);
	nand (gm_n377, gm_n88, in_24, gm_n76, gm_n376, gm_n141);
	nor (gm_n378, gm_n226, gm_n248, gm_n83, gm_n377);
	nand (gm_n379, gm_n361, gm_n144, gm_n124);
	nor (gm_n380, gm_n249, in_16, in_12, gm_n379, gm_n92);
	nand (gm_n381, gm_n141, in_24, in_20, gm_n380, gm_n205);
	nor (gm_n382, gm_n262, gm_n138, gm_n83, gm_n381);
	or (gm_n383, in_7, in_6, in_5);
	or (gm_n384, gm_n383, gm_n271);
	nor (gm_n385, gm_n188, gm_n63, in_8, gm_n384, gm_n282);
	nand (gm_n386, gm_n90, gm_n76, in_16, gm_n385, gm_n103);
	nor (gm_n387, gm_n214, gm_n83, gm_n82, gm_n386, gm_n216);
	nor (gm_n388, gm_n387, gm_n382, gm_n378);
	nand (gm_n389, gm_n351, gm_n172, gm_n163, gm_n388, gm_n373);
	nor (gm_n390, gm_n100, in_29, gm_n83);
	nor (gm_n391, in_26, in_25, gm_n82);
	and (gm_n392, in_18, in_17, in_16);
	not (gm_n393, gm_n392);
	nor (gm_n394, gm_n66, in_9, gm_n124);
	not (gm_n395, gm_n394);
	nor (gm_n396, in_2, in_1, gm_n94, in_4, in_3);
	nand (gm_n397, gm_n396, gm_n218);
	nand (gm_n398, gm_n64, gm_n175, in_12);
	or (gm_n399, gm_n395, gm_n62, gm_n61, gm_n398, gm_n397);
	nor (gm_n400, gm_n297, gm_n158, gm_n58, gm_n399, gm_n393);
	nand (gm_n401, gm_n390, in_31, gm_n54, gm_n400, gm_n391);
	nor (gm_n402, in_2, gm_n67, gm_n94, gm_n113, in_3);
	and (gm_n403, gm_n167, gm_n63, in_8, gm_n402, gm_n310);
	nor (gm_n404, in_16, gm_n62, in_14);
	nor (gm_n405, in_20, in_19, gm_n106);
	and (gm_n406, gm_n403, in_17, gm_n175, gm_n405, gm_n404);
	nor (gm_n407, in_24, in_23, in_22);
	nor (gm_n408, gm_n83, in_27, gm_n59);
	and (gm_n409, gm_n406, gm_n133, in_21, gm_n408, gm_n407);
	nand (gm_n410, gm_n55, gm_n100, in_29, gm_n409);
	not (gm_n411, gm_n255);
	not (gm_n412, gm_n270);
	nand (gm_n413, gm_n218, gm_n69, gm_n124);
	or (gm_n414, gm_n249, gm_n73, gm_n63, gm_n413, gm_n352);
	nor (gm_n415, gm_n411, gm_n82, gm_n76, gm_n414, gm_n412);
	nand (gm_n416, gm_n367, gm_n137, gm_n83, gm_n415);
	nand (gm_n417, gm_n416, gm_n410, gm_n401);
	and (gm_n418, gm_n310, gm_n208, gm_n124);
	nand (gm_n419, gm_n91, in_16, in_12, gm_n418, gm_n167);
	nor (gm_n420, gm_n165, gm_n82, gm_n76, gm_n419, gm_n206);
	nand (gm_n421, gm_n102, gm_n81, in_28, gm_n420);
	not (gm_n422, gm_n309);
	not (gm_n423, gm_n390);
	nor (gm_n424, in_10, in_9, in_8);
	nand (gm_n425, in_14, in_13, gm_n63);
	not (gm_n426, gm_n425);
	and (gm_n427, gm_n264, gm_n208, gm_n61, gm_n426, gm_n424);
	nand (gm_n428, gm_n173, in_19, in_15, gm_n427, gm_n359);
	nor (gm_n429, gm_n422, in_27, gm_n158, gm_n428, gm_n423);
	nand (gm_n430, gm_n429, in_31);
	not (gm_n431, gm_n358);
	not (gm_n432, gm_n65);
	nand (gm_n433, gm_n66, in_9, gm_n124);
	nand (gm_n434, in_6, gm_n70, in_4, gm_n320, in_7);
	or (gm_n435, gm_n432, in_15, gm_n61, gm_n434, gm_n433);
	nor (gm_n436, gm_n431, gm_n158, gm_n58, gm_n435, gm_n393);
	nand (gm_n437, gm_n100, in_29, in_28);
	not (gm_n438, gm_n437);
	nand (gm_n439, gm_n391, in_31, in_27, gm_n438, gm_n436);
	nand (gm_n440, gm_n439, gm_n430, gm_n421);
	nor (gm_n441, gm_n389, gm_n149, gm_n136, gm_n440, gm_n417);
	nand (gm_n442, gm_n110, gm_n63, in_8, gm_n208, gm_n189);
	nor (gm_n443, gm_n197, in_20, in_16, gm_n442, gm_n374);
	nand (gm_n444, gm_n103, in_28, in_24, gm_n443, gm_n367);
	nor (gm_n445, gm_n444, gm_n214);
	nor (gm_n446, in_15, gm_n64, gm_n175);
	nand (gm_n447, gm_n151, in_6, gm_n70);
	nor (gm_n448, gm_n447, gm_n114, in_8);
	and (gm_n449, gm_n446, gm_n73, in_12, gm_n448, gm_n228);
	nand (gm_n450, gm_n103, gm_n82, gm_n76, gm_n449, gm_n107);
	nor (gm_n451, gm_n216, gm_n195, gm_n83, gm_n450);
	not (gm_n452, gm_n173);
	nor (gm_n453, in_2, gm_n67, gm_n94, in_4, gm_n68);
	nand (gm_n454, gm_n189, gm_n65, in_11, gm_n453, gm_n394);
	nor (gm_n455, gm_n106, gm_n105, in_16);
	not (gm_n456, gm_n455);
	nor (gm_n457, gm_n452, gm_n58, in_15, gm_n456, gm_n454);
	nand (gm_n458, in_26, in_25, in_24);
	not (gm_n459, gm_n458);
	nand (gm_n460, gm_n308, in_27, in_23, gm_n459, gm_n457);
	nor (gm_n461, gm_n460, in_31);
	nor (gm_n462, gm_n461, gm_n451, gm_n445);
	not (gm_n463, gm_n235);
	nand (gm_n464, gm_n256, in_12, in_8, gm_n402, gm_n310);
	nor (gm_n465, gm_n236, gm_n76, in_16, gm_n464, gm_n463);
	nor (gm_n466, gm_n54, in_26, gm_n133);
	nand (gm_n467, gm_n227, in_28, in_24, gm_n466, gm_n465);
	nor (gm_n468, gm_n467, gm_n226);
	nand (gm_n469, in_2, in_1, in_0, in_4, in_3);
	nor (gm_n470, gm_n151, gm_n115, gm_n70, gm_n469, in_8);
	and (gm_n471, gm_n142, gm_n73, in_12, gm_n470, gm_n167);
	nand (gm_n472, gm_n107, gm_n82, in_20, gm_n471, gm_n263);
	nor (gm_n473, gm_n368, gm_n226, gm_n83, gm_n472);
	nand (gm_n474, gm_n310, gm_n257, gm_n124);
	nor (gm_n475, gm_n143, gm_n73, gm_n63, gm_n474, gm_n154);
	nand (gm_n476, gm_n58, gm_n106, in_17);
	not (gm_n477, gm_n476);
	nand (gm_n478, gm_n103, gm_n82, gm_n76, gm_n477, gm_n475);
	nand (gm_n479, gm_n55, in_30, in_29);
	nor (gm_n480, gm_n478, gm_n140, in_28, gm_n479);
	nor (gm_n481, gm_n480, gm_n473, gm_n468);
	nand (gm_n482, gm_n441, gm_n120, gm_n99, gm_n481, gm_n462);
	nand (gm_n483, gm_n70, gm_n113, gm_n68, gm_n145, gm_n115);
	nor (gm_n484, in_9, gm_n124, in_7, gm_n483, gm_n66);
	and (gm_n485, in_13, in_12);
	nor (gm_n486, gm_n105, gm_n73, in_15);
	nand (gm_n487, gm_n484, in_14, in_11, gm_n486, gm_n485);
	nor (gm_n488, in_21, in_20, in_19);
	not (gm_n489, gm_n488);
	nand (gm_n490, gm_n133, in_24, gm_n158);
	nor (gm_n491, gm_n487, in_22, in_18, gm_n490, gm_n489);
	nor (gm_n492, gm_n80, in_28, in_27);
	nand (gm_n493, in_31, gm_n100, gm_n59, gm_n492, gm_n491);
	nand (gm_n494, gm_n166, gm_n73, gm_n63, gm_n418, gm_n340);
	nor (gm_n495, gm_n206, gm_n82, gm_n76, gm_n494, gm_n412);
	and (gm_n496, in_31, in_30, in_29);
	nand (gm_n497, gm_n495, gm_n215, gm_n83, gm_n496);
	or (gm_n498, gm_n236, in_16, in_12, gm_n290, gm_n282);
	nor (gm_n499, gm_n206, gm_n82, in_20, gm_n498, gm_n412);
	nand (gm_n500, gm_n215, gm_n101, in_28, gm_n499);
	nand (gm_n501, gm_n500, gm_n497, gm_n493);
	nor (gm_n502, in_2, in_1, gm_n94, gm_n113, in_3);
	nand (gm_n503, gm_n502, gm_n144);
	nor (gm_n504, gm_n109, gm_n63, in_8, gm_n503, gm_n282);
	nand (gm_n505, gm_n90, in_20, in_16, gm_n504, gm_n227);
	nor (gm_n506, gm_n214, in_28, in_24, gm_n505, gm_n368);
	nor (out_0, gm_n501, gm_n482, gm_n79, gm_n506);
	and (gm_n508, gm_n150, gm_n73, gm_n63, gm_n448, gm_n167);
	nand (gm_n509, gm_n88, in_24, gm_n76, gm_n508, gm_n164);
	nor (gm_n510, gm_n226, gm_n216, gm_n83, gm_n509);
	nor (gm_n511, in_30, gm_n80, in_28);
	not (gm_n512, gm_n60);
	nor (gm_n513, gm_n87, in_21, in_20);
	not (gm_n514, gm_n513);
	nor (gm_n515, in_7, gm_n115, gm_n70);
	and (gm_n516, gm_n515, gm_n219, gm_n124);
	nand (gm_n517, gm_n302, gm_n340, in_15, gm_n516, gm_n426);
	nor (gm_n518, gm_n512, gm_n158, in_19, gm_n517, gm_n514);
	nand (gm_n519, gm_n511, in_31, in_27, gm_n518);
	not (gm_n520, gm_n227);
	and (gm_n521, in_19, in_18, in_17);
	not (gm_n522, gm_n521);
	nor (gm_n523, gm_n229, gm_n93);
	nand (gm_n524, gm_n142, gm_n63, gm_n124, gm_n523, gm_n340);
	nor (gm_n525, gm_n520, gm_n76, gm_n73, gm_n524, gm_n522);
	nand (gm_n526, gm_n81, in_28, gm_n82, gm_n525, gm_n215);
	nand (gm_n527, gm_n208, gm_n71, gm_n124);
	nor (gm_n528, gm_n236, gm_n73, in_12, gm_n527, gm_n288);
	nand (gm_n529, gm_n141, in_24, gm_n76, gm_n528, gm_n205);
	nor (gm_n530, gm_n216, gm_n234, gm_n83, gm_n529);
	nor (gm_n531, gm_n76, in_19, gm_n106);
	not (gm_n532, gm_n531);
	and (gm_n533, in_16, in_15, in_14);
	not (gm_n534, gm_n533);
	nand (gm_n535, in_5, gm_n113, gm_n68, gm_n145, gm_n115);
	nand (gm_n536, gm_n63, in_11, in_10);
	or (gm_n537, in_9, gm_n124, gm_n151, gm_n536, gm_n535);
	nor (gm_n538, gm_n532, gm_n105, in_13, gm_n537, gm_n534);
	nor (gm_n539, gm_n82, in_23, gm_n87);
	nor (gm_n540, in_28, gm_n54, in_26);
	nand (gm_n541, gm_n538, gm_n133, in_21, gm_n540, gm_n539);
	nor (gm_n542, gm_n55, in_30, gm_n80, gm_n541);
	and (gm_n543, in_2, in_1, in_0, in_3);
	and (gm_n544, gm_n115, in_5, gm_n113, gm_n543, gm_n151);
	nand (gm_n545, gm_n123, in_15, in_11, gm_n544, gm_n300);
	nor (gm_n546, gm_n393, in_23, in_19, gm_n545, gm_n514);
	nand (gm_n547, gm_n308, gm_n55, gm_n54, gm_n546, gm_n459);
	nand (gm_n548, in_2, gm_n67, in_0, gm_n113, gm_n68);
	nor (gm_n549, gm_n548, gm_n116, in_8);
	nand (gm_n550, gm_n110, gm_n73, in_12, gm_n549, gm_n207);
	nor (gm_n551, gm_n89, gm_n82, gm_n76, gm_n550, gm_n108);
	nand (gm_n552, gm_n225, gm_n139, gm_n83, gm_n551);
	nand (gm_n553, in_15, in_14, gm_n175);
	or (gm_n554, gm_n383, gm_n95);
	nor (gm_n555, gm_n553, gm_n63, in_8, gm_n554, gm_n282);
	nand (gm_n556, gm_n255, gm_n76, gm_n73, gm_n555, gm_n521);
	nor (gm_n557, gm_n234, gm_n83, gm_n82, gm_n556, gm_n85);
	nand (gm_n558, gm_n189, gm_n69, gm_n124);
	nor (gm_n559, gm_n109, gm_n73, in_12, gm_n558, gm_n237);
	nand (gm_n560, gm_n255, gm_n82, gm_n76, gm_n559, gm_n270);
	nor (gm_n561, gm_n224, gm_n185, in_28, gm_n560);
	nor (gm_n562, gm_n151, gm_n115, gm_n70, gm_n95, in_8);
	nand (gm_n563, gm_n200, in_16, in_12, gm_n562, gm_n256);
	nor (gm_n564, gm_n89, in_24, gm_n76, gm_n563, gm_n197);
	nand (gm_n565, gm_n496, gm_n139, gm_n83, gm_n564);
	not (gm_n566, gm_n217);
	nor (gm_n567, gm_n168, gm_n447, in_8);
	nand (gm_n568, gm_n153, in_16, gm_n63, gm_n567, gm_n207);
	nor (gm_n569, gm_n197, gm_n82, in_20, gm_n568, gm_n566);
	nand (gm_n570, gm_n496, gm_n84, in_28, gm_n569);
	nand (gm_n571, gm_n112, gm_n67, in_0, gm_n113, in_3);
	nor (gm_n572, gm_n571, gm_n345, gm_n124);
	and (gm_n573, gm_n150, in_16, gm_n63, gm_n572, gm_n242);
	nand (gm_n574, gm_n141, in_24, in_20, gm_n573, gm_n255);
	nor (gm_n575, gm_n479, gm_n262, gm_n83, gm_n574);
	and (gm_n576, gm_n199, in_16, in_12, gm_n346, gm_n150);
	nand (gm_n577, gm_n141, gm_n82, in_20, gm_n576, gm_n255);
	nor (gm_n578, gm_n368, gm_n234, gm_n83, gm_n577);
	nand (gm_n579, gm_n228, gm_n128, in_8, gm_n310);
	nor (gm_n580, gm_n314, in_19, gm_n62, gm_n579, gm_n456);
	nand (gm_n581, gm_n134, gm_n54, in_23, gm_n580, gm_n316);
	nor (gm_n582, gm_n581, gm_n423, gm_n55);
	not (gm_n583, gm_n391);
	nand (gm_n584, in_6, in_5, gm_n113, gm_n543, in_7);
	nor (gm_n585, gm_n395, in_15, in_11, gm_n584, gm_n398);
	nand (gm_n586, gm_n121, gm_n158, in_19, gm_n585, gm_n130);
	nor (gm_n587, gm_n357, gm_n55, gm_n54, gm_n586, gm_n583);
	nor (gm_n588, gm_n112, in_1, gm_n94, in_4, gm_n68);
	and (gm_n589, gm_n588, gm_n310, gm_n124);
	and (gm_n590, gm_n142, in_16, in_12, gm_n589, gm_n242);
	nand (gm_n591, gm_n90, gm_n82, in_20, gm_n590, gm_n103);
	nor (gm_n592, gm_n185, gm_n85, gm_n83, gm_n591);
	nor (gm_n593, gm_n582, gm_n578, gm_n575, gm_n592, gm_n587);
	nor (gm_n594, gm_n112, gm_n67, in_0, in_4, gm_n68);
	and (gm_n595, gm_n594, gm_n127, in_8);
	and (gm_n596, gm_n153, gm_n73, gm_n63, gm_n595, gm_n207);
	nand (gm_n597, gm_n141, gm_n82, gm_n76, gm_n596, gm_n205);
	nor (gm_n598, gm_n226, gm_n216, gm_n83, gm_n597);
	not (gm_n599, gm_n167);
	or (gm_n600, gm_n151, gm_n115, gm_n70, gm_n271);
	nor (gm_n601, gm_n599, in_12, gm_n124, gm_n600, gm_n177);
	nand (gm_n602, gm_n164, gm_n76, gm_n73, gm_n601, gm_n192);
	nor (gm_n603, gm_n224, in_28, gm_n82, gm_n602, gm_n214);
	nand (gm_n604, gm_n218, gm_n63, in_8, gm_n311, gm_n110);
	nor (gm_n605, gm_n553, in_20, gm_n73, gm_n604, gm_n476);
	nand (gm_n606, gm_n255, in_28, in_24, gm_n605, gm_n339);
	nor (gm_n607, gm_n606, gm_n185);
	nor (gm_n608, gm_n607, gm_n603, gm_n598);
	nor (gm_n609, gm_n92, gm_n73, in_12, gm_n266, gm_n553);
	nand (gm_n610, gm_n164, gm_n82, in_20, gm_n609, gm_n263);
	nor (gm_n611, gm_n262, gm_n226, in_28, gm_n610);
	not (gm_n612, gm_n337);
	nand (gm_n613, gm_n106, in_17, in_16);
	or (gm_n614, gm_n229, gm_n92, in_8, gm_n345);
	nor (gm_n615, gm_n432, gm_n58, in_15, gm_n614, gm_n613);
	nand (gm_n616, gm_n296, gm_n54, in_23, gm_n615, gm_n309);
	nor (gm_n617, gm_n616, gm_n612, in_31);
	not (gm_n618, gm_n306);
	not (gm_n619, gm_n424);
	nor (gm_n620, in_2, in_1, gm_n94, gm_n113, gm_n68);
	nand (gm_n621, gm_n620, gm_n218);
	nor (gm_n622, in_14, in_13, in_12);
	not (gm_n623, gm_n622);
	nor (gm_n624, gm_n619, in_15, in_11, gm_n623, gm_n621);
	nand (gm_n625, gm_n74, gm_n158, gm_n58, gm_n624, gm_n173);
	nor (gm_n626, gm_n618, in_31, gm_n54, gm_n625, gm_n422);
	nor (gm_n627, gm_n626, gm_n617, gm_n611);
	nand (gm_n628, gm_n593, gm_n570, gm_n565, gm_n627, gm_n608);
	not (gm_n629, gm_n479);
	not (gm_n630, gm_n263);
	or (gm_n631, gm_n345, gm_n95, in_8);
	or (gm_n632, gm_n188, gm_n73, in_12, gm_n631, gm_n352);
	nor (gm_n633, gm_n630, in_24, gm_n76, gm_n632, gm_n412);
	nand (gm_n634, gm_n629, gm_n367, in_28, gm_n633);
	nor (gm_n635, gm_n198, gm_n124, in_7, gm_n535, in_10);
	nor (gm_n636, gm_n175, in_12, in_11);
	nand (gm_n637, gm_n486, gm_n106, gm_n64, gm_n636, gm_n635);
	nand (gm_n638, gm_n86, in_20, in_19);
	nor (gm_n639, gm_n133, in_24, gm_n158);
	not (gm_n640, gm_n639);
	nor (gm_n641, gm_n637, in_26, gm_n87, gm_n640, gm_n638);
	nor (gm_n642, gm_n80, gm_n83, in_27);
	nand (gm_n643, gm_n641, gm_n55, in_30, gm_n642);
	and (gm_n644, gm_n199, gm_n63, gm_n124, gm_n402, gm_n218);
	nand (gm_n645, gm_n90, gm_n76, gm_n73, gm_n644, gm_n91);
	nor (gm_n646, gm_n104, gm_n83, gm_n82, gm_n645, gm_n216);
	nand (gm_n647, gm_n646, gm_n81);
	nand (gm_n648, gm_n647, gm_n643, gm_n634);
	nor (gm_n649, gm_n447, gm_n63, in_8, gm_n352, gm_n178);
	and (gm_n650, gm_n531, in_17, in_13, gm_n649, gm_n533);
	nor (gm_n651, in_24, gm_n158, gm_n87);
	and (gm_n652, gm_n408, in_25, gm_n86, gm_n651, gm_n650);
	nand (gm_n653, gm_n55, in_30, gm_n80, gm_n652);
	nand (gm_n654, gm_n208, gm_n189, gm_n124);
	nor (gm_n655, gm_n237, gm_n143, in_12, gm_n654);
	and (gm_n656, gm_n121, gm_n158, in_19, gm_n655, gm_n334);
	nor (gm_n657, in_26, gm_n133, in_24);
	nand (gm_n658, gm_n511, in_31, in_27, gm_n657, gm_n656);
	nand (gm_n659, gm_n150, in_16, gm_n63, gm_n595, gm_n242);
	nor (gm_n660, gm_n630, in_24, in_20, gm_n659, gm_n412);
	nand (gm_n661, gm_n186, gm_n137, gm_n83, gm_n660);
	nand (gm_n662, gm_n661, gm_n658, gm_n653);
	nor (gm_n663, gm_n628, gm_n561, gm_n557, gm_n662, gm_n648);
	nand (gm_n664, in_10, in_9, in_8);
	or (gm_n665, gm_n363, gm_n93, in_11, gm_n664, gm_n571);
	nor (gm_n666, gm_n514, gm_n58, gm_n62, gm_n665, gm_n613);
	nand (gm_n667, gm_n56, gm_n54, gm_n158, gm_n666, gm_n391);
	nor (gm_n668, gm_n667, gm_n55);
	nand (gm_n669, in_14, gm_n175, gm_n63);
	nand (gm_n670, in_10, gm_n198, gm_n124);
	nand (gm_n671, in_6, in_5, gm_n113, gm_n543, gm_n151);
	nor (gm_n672, gm_n669, in_15, in_11, gm_n671, gm_n670);
	nand (gm_n673, gm_n77, in_23, gm_n58, gm_n672, gm_n392);
	nor (gm_n674, in_30, in_29, gm_n83);
	not (gm_n675, gm_n674);
	nor (gm_n676, gm_n458, in_31, in_27, gm_n675, gm_n673);
	nor (gm_n677, gm_n322, in_15, gm_n61, gm_n434, gm_n363);
	nand (gm_n678, gm_n296, gm_n158, gm_n58, gm_n677, gm_n455);
	nor (gm_n679, gm_n57, gm_n55, in_27, gm_n678, gm_n422);
	nor (gm_n680, gm_n679, gm_n676, gm_n668);
	nor (gm_n681, gm_n92, in_16, gm_n63, gm_n290, gm_n374);
	nand (gm_n682, gm_n192, in_24, gm_n76, gm_n681, gm_n270);
	nor (gm_n683, gm_n216, gm_n195, in_28, gm_n682);
	not (gm_n684, gm_n496);
	and (gm_n685, gm_n320, in_8, in_4, gm_n515);
	and (gm_n686, gm_n153, in_16, gm_n63, gm_n685, gm_n446);
	nand (gm_n687, gm_n88, gm_n82, in_20, gm_n686, gm_n270);
	nor (gm_n688, gm_n684, gm_n368, gm_n83, gm_n687);
	nand (gm_n689, gm_n453, gm_n310, gm_n124);
	nor (gm_n690, gm_n109, in_16, gm_n63, gm_n689, gm_n154);
	nand (gm_n691, gm_n205, in_24, in_20, gm_n690, gm_n521);
	nor (gm_n692, gm_n138, gm_n224, in_28, gm_n691);
	nor (gm_n693, gm_n692, gm_n688, gm_n683);
	nand (gm_n694, gm_n663, gm_n552, gm_n547, gm_n693, gm_n680);
	nand (gm_n695, gm_n176, gm_n73, gm_n63, gm_n685, gm_n228);
	nor (gm_n696, gm_n165, in_24, gm_n76, gm_n695, gm_n411);
	nand (gm_n697, gm_n339, gm_n225, in_28, gm_n696);
	not (gm_n698, gm_n363);
	nor (gm_n699, gm_n277, gm_n447);
	nand (gm_n700, gm_n300, in_15, in_11, gm_n699, gm_n698);
	nor (gm_n701, gm_n317, in_23, in_19, gm_n700, gm_n456);
	nand (gm_n702, gm_n182, gm_n55, gm_n54, gm_n701, gm_n337);
	nor (gm_n703, in_2, gm_n67, in_0, gm_n113, gm_n68);
	and (gm_n704, gm_n703, gm_n144, in_8);
	nand (gm_n705, gm_n91, gm_n73, in_12, gm_n704, gm_n256);
	nor (gm_n706, gm_n206, gm_n82, in_20, gm_n705, gm_n463);
	nand (gm_n707, gm_n496, gm_n339, in_28, gm_n706);
	nand (gm_n708, gm_n707, gm_n702, gm_n697);
	nor (gm_n709, gm_n229, gm_n152, in_8);
	nand (gm_n710, gm_n142, in_16, in_12, gm_n709, gm_n340);
	nor (gm_n711, gm_n566, gm_n82, in_20, gm_n710, gm_n463);
	nand (gm_n712, gm_n139, gm_n81, in_28, gm_n711);
	nor (gm_n713, gm_n152, in_12, in_8, gm_n548, gm_n282);
	nand (gm_n714, gm_n200, in_20, in_16, gm_n713, gm_n164);
	nor (gm_n715, gm_n411, in_28, gm_n82, gm_n714, gm_n368);
	nand (gm_n716, gm_n715, gm_n496);
	or (gm_n717, gm_n143, gm_n73, in_12, gm_n689, gm_n237);
	nor (gm_n718, gm_n165, in_24, gm_n76, gm_n717, gm_n206);
	nand (gm_n719, gm_n496, gm_n139, in_28, gm_n718);
	nand (gm_n720, gm_n719, gm_n716, gm_n712);
	nor (gm_n721, gm_n694, gm_n542, gm_n530, gm_n720, gm_n708);
	nor (gm_n722, gm_n109, in_16, gm_n63, gm_n290, gm_n111);
	nand (gm_n723, gm_n192, gm_n82, in_20, gm_n722, gm_n270);
	nor (gm_n724, gm_n479, gm_n224, gm_n83, gm_n723);
	nand (gm_n725, gm_n66, in_9, in_8);
	nand (gm_n726, gm_n208, gm_n127);
	nor (gm_n727, gm_n725, in_15, in_11, gm_n726, gm_n669);
	nand (gm_n728, gm_n121, gm_n158, in_19, gm_n727, gm_n513);
	nor (gm_n729, gm_n183, gm_n55, gm_n54, gm_n728, gm_n612);
	and (gm_n730, in_10, in_9, in_8);
	nor (gm_n731, gm_n112, in_1, in_0, in_4, in_3);
	and (gm_n732, gm_n144, gm_n175, in_11, gm_n731, gm_n730);
	nor (gm_n733, gm_n73, gm_n62, in_14);
	and (gm_n734, gm_n405, in_17, in_12, gm_n733, gm_n732);
	nor (gm_n735, gm_n83, in_27, in_26);
	nand (gm_n736, gm_n407, in_25, in_21, gm_n735, gm_n734);
	nor (gm_n737, in_31, gm_n100, in_29, gm_n736);
	nor (gm_n738, gm_n737, gm_n729, gm_n724);
	nand (gm_n739, gm_n144, gm_n128);
	nor (gm_n740, gm_n236, gm_n63, gm_n124, gm_n739, gm_n237);
	nand (gm_n741, gm_n192, in_20, in_16, gm_n740, gm_n521);
	nor (gm_n742, gm_n138, in_28, in_24, gm_n741, gm_n368);
	nand (gm_n743, gm_n110, gm_n63, gm_n124, gm_n731, gm_n264);
	nor (gm_n744, gm_n187, in_20, gm_n73, gm_n743, gm_n143);
	nand (gm_n745, gm_n339, in_28, gm_n82, gm_n744, gm_n263);
	nor (gm_n746, gm_n745, gm_n226);
	nand (gm_n747, gm_n66, in_9, gm_n124, gm_n310, gm_n219);
	nor (gm_n748, gm_n122, gm_n62, gm_n61, gm_n747, gm_n669);
	nand (gm_n749, gm_n60, in_23, gm_n58, gm_n748, gm_n130);
	nor (gm_n750, gm_n612, gm_n55, gm_n54, gm_n749);
	nor (gm_n751, gm_n750, gm_n746, gm_n742);
	nand (gm_n752, gm_n721, gm_n526, gm_n519, gm_n751, gm_n738);
	nand (gm_n753, gm_n112, in_1, in_0, gm_n113, in_3);
	nor (gm_n754, gm_n753, gm_n116, in_8);
	nand (gm_n755, gm_n150, gm_n73, gm_n63, gm_n754, gm_n153);
	nor (gm_n756, gm_n463, in_24, gm_n76, gm_n755, gm_n411);
	nand (gm_n757, gm_n213, gm_n139, gm_n83, gm_n756);
	nand (gm_n758, gm_n115, gm_n70, in_4, gm_n320, gm_n151);
	or (gm_n759, gm_n432, in_15, gm_n61, gm_n758, gm_n725);
	nor (gm_n760, gm_n452, in_23, in_19, gm_n759, gm_n303);
	nand (gm_n761, gm_n134, in_31, in_27, gm_n760, gm_n390);
	or (gm_n762, gm_n177, gm_n73, in_12, gm_n282, gm_n238);
	nor (gm_n763, gm_n104, gm_n82, gm_n76, gm_n762, gm_n108);
	nand (gm_n764, gm_n466, gm_n196, gm_n83, gm_n763);
	nand (gm_n765, gm_n764, gm_n761, gm_n757);
	or (gm_n766, gm_n152, gm_n63, gm_n124, gm_n352, gm_n95);
	nand (gm_n767, in_16, gm_n62, gm_n64);
	nor (gm_n768, gm_n157, gm_n105, gm_n175, gm_n767, gm_n766);
	nor (gm_n769, in_24, in_23, gm_n87);
	and (gm_n770, in_28, in_27, in_26);
	nand (gm_n771, gm_n768, in_25, in_21, gm_n770, gm_n769);
	nor (gm_n772, gm_n55, gm_n100, gm_n80, gm_n771);
	nor (out_1, gm_n765, gm_n752, gm_n510, gm_n772);
	not (gm_n774, gm_n466);
	nor (gm_n775, gm_n112, in_1, gm_n94, in_4, in_3);
	nand (gm_n776, gm_n775, gm_n189, in_8);
	nor (gm_n777, gm_n92, in_16, gm_n63, gm_n776, gm_n188);
	nand (gm_n778, gm_n90, gm_n82, in_20, gm_n777, gm_n192);
	nor (gm_n779, gm_n774, gm_n195, gm_n83, gm_n778);
	nor (gm_n780, gm_n152, gm_n63, gm_n124, gm_n168, gm_n111);
	nand (gm_n781, gm_n164, gm_n76, in_16, gm_n780, gm_n166);
	nor (gm_n782, gm_n248, in_28, in_24, gm_n781, gm_n520);
	nand (gm_n783, gm_n782, gm_n213);
	nor (gm_n784, gm_n271, gm_n447, gm_n124);
	nand (gm_n785, gm_n91, in_16, gm_n63, gm_n784, gm_n256);
	nor (gm_n786, gm_n89, gm_n82, gm_n76, gm_n785, gm_n522);
	nand (gm_n787, gm_n213, gm_n186, gm_n83, gm_n786);
	nand (gm_n788, gm_n144, in_12, gm_n124, gm_n703, gm_n153);
	nor (gm_n789, gm_n165, in_20, in_16, gm_n788, gm_n188);
	nand (gm_n790, gm_n255, in_28, gm_n82, gm_n789, gm_n339);
	nor (gm_n791, gm_n790, gm_n214);
	and (gm_n792, in_6, gm_n70, gm_n113, gm_n543, in_7);
	and (gm_n793, gm_n426, gm_n62, gm_n61, gm_n792, gm_n730);
	nand (gm_n794, gm_n316, in_23, in_19, gm_n793, gm_n359);
	nor (gm_n795, gm_n183, in_31, in_27, gm_n794, gm_n612);
	not (gm_n796, gm_n74);
	not (gm_n797, gm_n725);
	nand (gm_n798, gm_n65, in_15, in_11, gm_n332, gm_n797);
	nor (gm_n799, gm_n796, gm_n158, in_19, gm_n798, gm_n335);
	nand (gm_n800, gm_n337, in_31, gm_n54, gm_n799, gm_n657);
	not (gm_n801, gm_n192);
	nand (gm_n802, gm_n176, gm_n73, gm_n63, gm_n341, gm_n256);
	nor (gm_n803, gm_n165, gm_n82, in_20, gm_n802, gm_n801);
	nand (gm_n804, gm_n367, gm_n196, gm_n83, gm_n803);
	nand (gm_n805, gm_n218, gm_n63, gm_n124, gm_n502, gm_n153);
	nor (gm_n806, gm_n108, gm_n76, in_16, gm_n805, gm_n143);
	nand (gm_n807, gm_n88, gm_n83, gm_n82, gm_n806, gm_n186);
	nor (gm_n808, gm_n807, gm_n195);
	nor (gm_n809, gm_n117, gm_n63, gm_n124, gm_n352, gm_n374);
	nand (gm_n810, gm_n235, gm_n76, gm_n73, gm_n809, gm_n255);
	nor (gm_n811, gm_n224, in_28, in_24, gm_n810, gm_n195);
	nand (gm_n812, gm_n446, gm_n76, gm_n73, gm_n270, gm_n209);
	nor (gm_n813, gm_n140, gm_n83, gm_n82, gm_n812, gm_n630);
	nand (gm_n814, gm_n813, gm_n213);
	nand (gm_n815, gm_n126, in_15, in_11, gm_n698, gm_n332);
	nor (gm_n816, gm_n796, in_23, in_19, gm_n815, gm_n317);
	nand (gm_n817, gm_n182, in_31, in_27, gm_n816, gm_n337);
	nand (gm_n818, gm_n199, gm_n63, gm_n124, gm_n257, gm_n189);
	nor (gm_n819, gm_n236, gm_n76, gm_n73, gm_n818, gm_n412);
	nand (gm_n820, gm_n88, in_28, gm_n82, gm_n819, gm_n339);
	nor (gm_n821, gm_n820, gm_n234);
	nand (gm_n822, gm_n264, gm_n128);
	nor (gm_n823, gm_n154, in_12, in_8, gm_n822, gm_n374);
	nand (gm_n824, gm_n192, gm_n76, in_16, gm_n823, gm_n235);
	nor (gm_n825, gm_n248, in_28, gm_n82, gm_n824, gm_n226);
	nor (gm_n826, gm_n725, gm_n62, gm_n61, gm_n758, gm_n314);
	nand (gm_n827, gm_n455, gm_n158, in_19, gm_n826, gm_n513);
	nor (gm_n828, gm_n512, in_31, gm_n54, gm_n827, gm_n437);
	nand (gm_n829, in_7, gm_n115, in_5, gm_n361, in_8);
	nor (gm_n830, gm_n109, in_16, in_12, gm_n829, gm_n599);
	nand (gm_n831, gm_n88, gm_n82, gm_n76, gm_n830, gm_n235);
	nor (gm_n832, gm_n85, gm_n234, in_28, gm_n831);
	or (gm_n833, gm_n447, in_12, in_8, gm_n271, gm_n282);
	nor (gm_n834, gm_n109, gm_n76, gm_n73, gm_n833, gm_n412);
	nand (gm_n835, gm_n103, gm_n83, gm_n82, gm_n834, gm_n139);
	nor (gm_n836, gm_n835, gm_n214);
	nor (gm_n837, gm_n828, gm_n825, gm_n821, gm_n836, gm_n832);
	not (gm_n838, gm_n511);
	nor (gm_n839, gm_n432, gm_n62, in_11, gm_n584, gm_n670);
	nand (gm_n840, gm_n316, in_23, in_19, gm_n839, gm_n392);
	nor (gm_n841, gm_n512, in_31, gm_n54, gm_n840, gm_n838);
	nand (gm_n842, gm_n515, gm_n69, in_8);
	nor (gm_n843, gm_n553, in_16, in_12, gm_n842, gm_n282);
	nand (gm_n844, gm_n217, gm_n82, gm_n76, gm_n843, gm_n235);
	nor (gm_n845, gm_n140, gm_n185, in_28, gm_n844);
	nor (gm_n846, in_9, gm_n124, gm_n151, gm_n483, gm_n66);
	nand (gm_n847, gm_n175, gm_n63, in_11, gm_n846, gm_n64);
	nor (gm_n848, in_17, in_16, gm_n62, gm_n847, in_18);
	and (gm_n849, gm_n488, in_26, in_22, gm_n848, gm_n639);
	and (gm_n850, gm_n642, gm_n55, gm_n100, gm_n849);
	nor (gm_n851, gm_n850, gm_n845, gm_n841);
	or (gm_n852, gm_n447, gm_n63, gm_n124, gm_n288, gm_n168);
	nor (gm_n853, gm_n188, gm_n76, in_16, gm_n852, gm_n412);
	nand (gm_n854, gm_n102, in_28, in_24, gm_n853, gm_n192);
	nor (gm_n855, gm_n854, gm_n234);
	nand (gm_n856, gm_n127, gm_n126, gm_n61, gm_n426, gm_n311);
	nor (gm_n857, gm_n796, in_19, gm_n62, gm_n856, gm_n297);
	nand (gm_n858, gm_n56, gm_n54, gm_n158, gm_n857, gm_n182);
	nor (gm_n859, gm_n858, in_31);
	or (gm_n860, gm_n152, in_12, gm_n124, gm_n229, gm_n92);
	nor (gm_n861, gm_n197, gm_n76, gm_n73, gm_n860, gm_n553);
	nand (gm_n862, gm_n103, gm_n83, in_24, gm_n861, gm_n139);
	nor (gm_n863, gm_n862, gm_n185);
	nor (gm_n864, gm_n863, gm_n859, gm_n855);
	nand (gm_n865, gm_n837, gm_n817, gm_n814, gm_n864, gm_n851);
	and (gm_n866, gm_n243, gm_n127, gm_n124);
	nand (gm_n867, gm_n166, in_16, in_12, gm_n866, gm_n242);
	nor (gm_n868, gm_n89, gm_n82, in_20, gm_n867, gm_n165);
	nand (gm_n869, gm_n102, gm_n81, in_28, gm_n868);
	nor (gm_n870, gm_n271, gm_n116, gm_n124);
	nand (gm_n871, gm_n91, gm_n73, in_12, gm_n870, gm_n167);
	nor (gm_n872, gm_n165, gm_n82, in_20, gm_n871, gm_n566);
	nand (gm_n873, gm_n225, gm_n84, in_28, gm_n872);
	nand (gm_n874, gm_n257, gm_n218);
	or (gm_n875, gm_n314, in_15, gm_n61, gm_n874, gm_n664);
	nor (gm_n876, gm_n122, gm_n158, in_19, gm_n875, gm_n297);
	nand (gm_n877, gm_n182, in_31, gm_n54, gm_n876, gm_n511);
	nand (gm_n878, gm_n877, gm_n873, gm_n869);
	and (gm_n879, gm_n775, gm_n144, in_8);
	nand (gm_n880, gm_n142, in_16, in_12, gm_n879, gm_n153);
	nor (gm_n881, gm_n463, in_24, gm_n76, gm_n880, gm_n630);
	nand (gm_n882, gm_n466, gm_n196, in_28, gm_n881);
	and (gm_n883, gm_n124, gm_n113, gm_n68, gm_n515, gm_n145);
	nand (gm_n884, gm_n167, in_16, gm_n63, gm_n883, gm_n446);
	nor (gm_n885, gm_n801, gm_n82, in_20, gm_n884, gm_n522);
	nand (gm_n886, gm_n196, gm_n84, gm_n83, gm_n885);
	nor (gm_n887, gm_n548, gm_n447, gm_n124);
	nand (gm_n888, gm_n166, in_16, gm_n63, gm_n887, gm_n340);
	nor (gm_n889, gm_n206, in_24, gm_n76, gm_n888, gm_n476);
	nand (gm_n890, gm_n629, gm_n84, in_28, gm_n889);
	nand (gm_n891, gm_n890, gm_n886, gm_n882);
	nor (gm_n892, gm_n865, gm_n811, gm_n808, gm_n891, gm_n878);
	nor (gm_n893, gm_n188, gm_n73, in_12, gm_n413, gm_n237);
	nand (gm_n894, gm_n88, in_24, gm_n76, gm_n893, gm_n164);
	nor (gm_n895, gm_n214, gm_n140, in_28, gm_n894);
	nand (gm_n896, gm_n311, gm_n218, gm_n124);
	nor (gm_n897, gm_n553, gm_n73, in_12, gm_n896, gm_n282);
	nand (gm_n898, gm_n227, in_24, in_20, gm_n897, gm_n521);
	nor (gm_n899, gm_n774, gm_n185, gm_n83, gm_n898);
	nor (gm_n900, gm_n571, gm_n116, gm_n124);
	and (gm_n901, gm_n199, in_16, in_12, gm_n900, gm_n150);
	nand (gm_n902, gm_n164, gm_n82, gm_n76, gm_n901, gm_n217);
	nor (gm_n903, gm_n684, gm_n368, in_28, gm_n902);
	nor (gm_n904, gm_n903, gm_n899, gm_n895);
	nand (gm_n905, gm_n243, gm_n218, in_8);
	nor (gm_n906, gm_n398, gm_n352, gm_n62, gm_n905, gm_n613);
	nand (gm_n907, gm_n309, in_23, gm_n58, gm_n906, gm_n513);
	nor (gm_n908, gm_n357, in_31, in_27, gm_n907);
	nand (gm_n909, gm_n620, gm_n71, gm_n124);
	nor (gm_n910, gm_n92, in_16, in_12, gm_n909, gm_n143);
	nand (gm_n911, gm_n205, in_24, in_20, gm_n910, gm_n521);
	nor (gm_n912, gm_n479, gm_n216, in_28, gm_n911);
	nor (gm_n913, gm_n345, gm_n271, gm_n124);
	and (gm_n914, gm_n446, in_16, gm_n63, gm_n913, gm_n242);
	nand (gm_n915, gm_n217, gm_n82, gm_n76, gm_n914, gm_n270);
	nor (gm_n916, gm_n262, gm_n195, gm_n83, gm_n915);
	nor (gm_n917, gm_n916, gm_n912, gm_n908);
	nand (gm_n918, gm_n892, gm_n804, gm_n800, gm_n917, gm_n904);
	nand (gm_n919, gm_n142, in_16, in_12, gm_n228, gm_n220);
	nor (gm_n920, gm_n566, in_24, in_20, gm_n919, gm_n522);
	nand (gm_n921, gm_n225, gm_n102, in_28, gm_n920);
	nor (gm_n922, gm_n188, in_16, gm_n63, gm_n474, gm_n288);
	and (gm_n923, gm_n103, in_24, in_20, gm_n922, gm_n521);
	nand (gm_n924, gm_n213, gm_n84, gm_n83, gm_n923);
	nand (gm_n925, gm_n394, gm_n189, gm_n61, gm_n453);
	or (gm_n926, gm_n432, in_19, gm_n62, gm_n925, gm_n393);
	nor (gm_n927, gm_n512, gm_n54, in_23, gm_n926, gm_n131);
	nand (gm_n928, gm_n927, gm_n511, gm_n55);
	nand (gm_n929, gm_n928, gm_n924, gm_n921);
	not (gm_n930, gm_n433);
	nor (gm_n931, in_14, in_13, gm_n63);
	nand (gm_n932, gm_n930, gm_n62, in_11, gm_n544, gm_n931);
	nor (gm_n933, gm_n297, in_23, in_19, gm_n932, gm_n456);
	nand (gm_n934, gm_n459, in_31, gm_n54, gm_n933, gm_n674);
	and (gm_n935, gm_n110, in_12, in_8, gm_n264, gm_n257);
	nand (gm_n936, gm_n142, gm_n76, in_16, gm_n935, gm_n235);
	nor (gm_n937, gm_n224, gm_n83, gm_n82, gm_n936, gm_n206);
	nand (gm_n938, gm_n937, gm_n137);
	or (gm_n939, gm_n352, gm_n796, gm_n62, gm_n905, gm_n623);
	nor (gm_n940, gm_n183, gm_n158, gm_n58, gm_n939, gm_n514);
	nand (gm_n941, gm_n308, gm_n55, gm_n54, gm_n940);
	nand (gm_n942, gm_n941, gm_n938, gm_n934);
	nor (gm_n943, gm_n918, gm_n795, gm_n791, gm_n942, gm_n929);
	or (gm_n944, gm_n151, gm_n115, gm_n70, gm_n95, gm_n124);
	nor (gm_n945, gm_n236, in_16, in_12, gm_n944, gm_n599);
	nand (gm_n946, gm_n227, gm_n82, gm_n76, gm_n945, gm_n235);
	nor (gm_n947, gm_n479, gm_n774, in_28, gm_n946);
	and (gm_n948, gm_n127, gm_n113, gm_n68, gm_n300, gm_n145);
	and (gm_n949, gm_n121, in_15, in_11, gm_n948, gm_n123);
	nand (gm_n950, gm_n316, in_23, in_19, gm_n949, gm_n657);
	nor (gm_n951, gm_n57, gm_n55, in_27, gm_n950);
	nand (gm_n952, gm_n402, gm_n189, in_8);
	nor (gm_n953, gm_n143, gm_n73, gm_n63, gm_n952, gm_n288);
	nand (gm_n954, gm_n90, gm_n82, gm_n76, gm_n953, gm_n192);
	nor (gm_n955, gm_n479, gm_n140, in_28, gm_n954);
	nor (gm_n956, gm_n955, gm_n951, gm_n947);
	nor (gm_n957, gm_n92, gm_n63, gm_n124, gm_n571, gm_n447);
	and (gm_n958, gm_n141, gm_n76, gm_n73, gm_n957, gm_n176);
	nand (gm_n959, gm_n84, gm_n83, in_24, gm_n958, gm_n88);
	nor (gm_n960, gm_n959, gm_n684);
	nor (gm_n961, gm_n345, gm_n178, gm_n124);
	and (gm_n962, gm_n446, gm_n73, gm_n63, gm_n961, gm_n228);
	nand (gm_n963, gm_n205, in_24, gm_n76, gm_n962, gm_n270);
	nor (gm_n964, gm_n138, gm_n85, gm_n83, gm_n963);
	nand (gm_n965, gm_n218, gm_n113, gm_n68, gm_n145);
	nor (gm_n966, gm_n111, gm_n63, gm_n124, gm_n965, gm_n374);
	nand (gm_n967, gm_n141, in_20, in_16, gm_n966, gm_n205);
	nor (gm_n968, gm_n368, in_28, in_24, gm_n967, gm_n684);
	nor (gm_n969, gm_n968, gm_n964, gm_n960);
	nand (gm_n970, gm_n943, gm_n787, gm_n783, gm_n969, gm_n956);
	nand (gm_n971, in_7, gm_n115, gm_n70);
	nand (gm_n972, gm_n112, gm_n67, gm_n94, in_4, in_3);
	nor (gm_n973, gm_n972, gm_n971);
	nand (gm_n974, gm_n142, in_12, gm_n124, gm_n973, gm_n256);
	nor (gm_n975, gm_n566, gm_n76, in_16, gm_n974, gm_n463);
	nand (gm_n976, gm_n84, in_28, gm_n82, gm_n975, gm_n496);
	not (gm_n977, gm_n657);
	or (gm_n978, gm_n669, gm_n62, in_11, gm_n393, gm_n362);
	nor (gm_n979, gm_n335, in_23, gm_n58, gm_n978, gm_n977);
	nand (gm_n980, gm_n390, gm_n55, in_27, gm_n979);
	and (gm_n981, gm_n124, in_4, gm_n68, gm_n145, gm_n144);
	nand (gm_n982, gm_n199, in_16, in_12, gm_n981, gm_n150);
	nor (gm_n983, gm_n801, gm_n82, in_20, gm_n982, gm_n522);
	nand (gm_n984, gm_n215, gm_n196, gm_n83, gm_n983);
	nand (gm_n985, gm_n984, gm_n980, gm_n976);
	nand (gm_n986, gm_n115, in_5, gm_n113, gm_n543, in_7);
	nor (gm_n987, gm_n363, in_15, gm_n61, gm_n986, gm_n619);
	nand (gm_n988, gm_n358, in_23, in_19, gm_n987, gm_n455);
	nor (gm_n989, gm_n618, in_31, in_27, gm_n988, gm_n583);
	nor (out_2, gm_n985, gm_n970, gm_n779, gm_n989);
	nand (gm_n991, gm_n64, in_13, gm_n63);
	nor (gm_n992, gm_n125, in_15, in_11, gm_n991, gm_n874);
	nand (gm_n993, gm_n121, in_23, gm_n58, gm_n992, gm_n296);
	nor (gm_n994, gm_n57, gm_n55, gm_n54, gm_n993, gm_n977);
	not (gm_n995, gm_n322);
	nand (gm_n996, gm_n289, gm_n264, in_11, gm_n995);
	or (gm_n997, gm_n363, gm_n58, in_15, gm_n996, gm_n613);
	nor (gm_n998, gm_n431, gm_n54, in_23, gm_n997, gm_n458);
	nand (gm_n999, gm_n998, gm_n511, gm_n55);
	and (gm_n1000, gm_n265, gm_n144);
	nand (gm_n1001, gm_n176, in_12, in_8, gm_n1000, gm_n228);
	nor (gm_n1002, gm_n165, gm_n76, gm_n73, gm_n1001, gm_n411);
	nand (gm_n1003, gm_n367, in_28, in_24, gm_n1002, gm_n629);
	nand (gm_n1004, gm_n167, in_12, in_8, gm_n264, gm_n243);
	nor (gm_n1005, gm_n108, in_20, in_16, gm_n1004, gm_n177);
	nand (gm_n1006, gm_n84, in_28, in_24, gm_n1005, gm_n255);
	nor (gm_n1007, gm_n1006, gm_n138);
	nor (gm_n1008, gm_n154, in_16, gm_n63, gm_n527, gm_n177);
	nand (gm_n1009, gm_n217, gm_n82, in_20, gm_n1008, gm_n235);
	nor (gm_n1010, gm_n214, gm_n248, gm_n83, gm_n1009);
	nor (gm_n1011, gm_n345, gm_n168, in_8);
	nand (gm_n1012, gm_n199, in_16, gm_n63, gm_n1011, gm_n150);
	nor (gm_n1013, gm_n108, in_24, gm_n76, gm_n1012, gm_n411);
	nand (gm_n1014, gm_n466, gm_n196, in_28, gm_n1013);
	nor (gm_n1015, gm_n271, gm_n971, gm_n124);
	nand (gm_n1016, gm_n153, in_16, in_12, gm_n1015, gm_n176);
	nor (gm_n1017, gm_n187, gm_n82, in_20, gm_n1016, gm_n566);
	nand (gm_n1018, gm_n225, gm_n84, gm_n83, gm_n1017);
	nand (gm_n1019, gm_n310, gm_n219, in_8);
	nor (gm_n1020, gm_n177, in_16, gm_n63, gm_n1019, gm_n237);
	nand (gm_n1021, gm_n217, gm_n82, gm_n76, gm_n1020, gm_n235);
	nor (gm_n1022, gm_n479, gm_n368, in_28, gm_n1021);
	or (gm_n1023, gm_n151, gm_n115, in_5, gm_n469, gm_n124);
	nor (gm_n1024, gm_n553, gm_n73, gm_n63, gm_n1023, gm_n599);
	nand (gm_n1025, gm_n263, in_24, gm_n76, gm_n1024, gm_n477);
	nor (gm_n1026, gm_n185, gm_n85, gm_n83, gm_n1025);
	or (gm_n1027, gm_n188, gm_n63, in_11, gm_n758, gm_n670);
	nor (gm_n1028, gm_n463, in_20, in_16, gm_n1027, gm_n411);
	nand (gm_n1029, gm_n84, in_28, in_24, gm_n1028, gm_n496);
	or (gm_n1030, gm_n321, gm_n62, gm_n61, gm_n425, gm_n322);
	nor (gm_n1031, gm_n122, gm_n158, gm_n58, gm_n1030, gm_n317);
	nand (gm_n1032, gm_n305, gm_n55, in_27, gm_n1031, gm_n438);
	not (gm_n1033, gm_n178);
	nand (gm_n1034, gm_n1033, gm_n144);
	nor (gm_n1035, gm_n92, in_12, gm_n124, gm_n1034, gm_n177);
	nand (gm_n1036, gm_n192, gm_n76, in_16, gm_n1035, gm_n270);
	nor (gm_n1037, gm_n216, gm_n83, in_24, gm_n1036, gm_n479);
	or (gm_n1038, gm_n383, gm_n178);
	nor (gm_n1039, gm_n322, in_15, gm_n61, gm_n1038, gm_n623);
	nand (gm_n1040, gm_n173, in_23, in_19, gm_n1039, gm_n359);
	nor (gm_n1041, gm_n618, gm_n55, in_27, gm_n1040, gm_n977);
	not (gm_n1042, gm_n613);
	nor (gm_n1043, gm_n670, gm_n62, in_11, gm_n600, gm_n363);
	nand (gm_n1044, gm_n513, in_23, in_19, gm_n1043, gm_n1042);
	nor (gm_n1045, gm_n422, gm_n55, in_27, gm_n1044, gm_n612);
	nand (gm_n1046, gm_n265, gm_n218, in_8);
	nor (gm_n1047, gm_n425, gm_n237, gm_n62, gm_n1046, gm_n456);
	nand (gm_n1048, gm_n459, gm_n158, gm_n58, gm_n1047, gm_n513);
	nor (gm_n1049, gm_n423, in_31, in_27, gm_n1048);
	nand (gm_n1050, in_28, in_27, gm_n59);
	nor (gm_n1051, gm_n73, gm_n62, in_14, gm_n323, gm_n105);
	nand (gm_n1052, gm_n326, in_25, in_21, gm_n1051, gm_n531);
	nor (gm_n1053, gm_n55, in_30, gm_n80, gm_n1052, gm_n1050);
	nor (gm_n1054, gm_n1045, gm_n1041, gm_n1037, gm_n1053, gm_n1049);
	nor (gm_n1055, gm_n971, gm_n95, gm_n124);
	and (gm_n1056, gm_n446, gm_n73, in_12, gm_n1055, gm_n340);
	nand (gm_n1057, gm_n90, gm_n82, gm_n76, gm_n1056, gm_n263);
	nor (gm_n1058, gm_n684, gm_n774, gm_n83, gm_n1057);
	or (gm_n1059, in_7, in_6, gm_n70, gm_n469, in_8);
	nor (gm_n1060, gm_n249, gm_n73, gm_n63, gm_n1059, gm_n599);
	nand (gm_n1061, gm_n88, in_24, in_20, gm_n1060, gm_n521);
	nor (gm_n1062, gm_n195, gm_n224, in_28, gm_n1061);
	or (gm_n1063, gm_n95, gm_n93, gm_n124);
	nor (gm_n1064, gm_n236, gm_n73, in_12, gm_n1063, gm_n282);
	nand (gm_n1065, gm_n90, in_24, in_20, gm_n1064, gm_n255);
	nor (gm_n1066, gm_n214, gm_n85, gm_n83, gm_n1065);
	nor (gm_n1067, gm_n1066, gm_n1062, gm_n1058);
	nand (gm_n1068, gm_n361, gm_n310, in_8);
	nor (gm_n1069, gm_n599, gm_n73, in_12, gm_n1068, gm_n374);
	nand (gm_n1070, gm_n263, gm_n82, in_20, gm_n1069, gm_n270);
	nor (gm_n1071, gm_n368, gm_n234, in_28, gm_n1070);
	nand (gm_n1072, gm_n167, in_12, gm_n124, gm_n502, gm_n515);
	nor (gm_n1073, gm_n108, gm_n76, gm_n73, gm_n1072, gm_n109);
	nand (gm_n1074, gm_n103, in_28, in_24, gm_n1073, gm_n466);
	nor (gm_n1075, gm_n1074, gm_n138);
	nor (gm_n1076, gm_n432, gm_n62, in_11, gm_n621, gm_n725);
	nand (gm_n1077, gm_n296, gm_n158, in_19, gm_n1076, gm_n359);
	nor (gm_n1078, gm_n357, in_31, gm_n54, gm_n1077, gm_n977);
	nor (gm_n1079, gm_n1078, gm_n1075, gm_n1071);
	nand (gm_n1080, gm_n1054, gm_n1032, gm_n1029, gm_n1079, gm_n1067);
	and (gm_n1081, gm_n115, in_5, in_4, gm_n320, in_7);
	nand (gm_n1082, gm_n65, gm_n62, in_11, gm_n1081, gm_n930);
	nor (gm_n1083, gm_n331, in_23, in_19, gm_n1082, gm_n297);
	nand (gm_n1084, gm_n390, in_31, in_27, gm_n1083, gm_n459);
	nand (gm_n1085, gm_n200, gm_n63, in_8, gm_n523, gm_n228);
	nor (gm_n1086, gm_n104, in_20, gm_n73, gm_n1085, gm_n108);
	nand (gm_n1087, gm_n139, gm_n83, gm_n82, gm_n1086, gm_n629);
	nand (gm_n1088, gm_n127, in_12, gm_n124, gm_n208, gm_n167);
	or (gm_n1089, gm_n249, in_20, gm_n73, gm_n1088, gm_n165);
	nor (gm_n1090, gm_n104, gm_n83, gm_n82, gm_n1089, gm_n774);
	nand (gm_n1091, gm_n1090, gm_n101);
	nand (gm_n1092, gm_n1091, gm_n1087, gm_n1084);
	nand (gm_n1093, gm_n153, gm_n73, gm_n63, gm_n278, gm_n176);
	nor (gm_n1094, gm_n566, gm_n82, gm_n76, gm_n1093, gm_n522);
	nand (gm_n1095, gm_n496, gm_n215, in_28, gm_n1094);
	nor (gm_n1096, gm_n670, gm_n447, in_11, gm_n753, gm_n398);
	nand (gm_n1097, gm_n296, gm_n58, gm_n62, gm_n1096, gm_n359);
	nor (gm_n1098, gm_n57, in_27, in_23, gm_n1097, gm_n458);
	nand (gm_n1099, gm_n1098, gm_n55);
	nand (gm_n1100, in_8, gm_n113, gm_n68, gm_n515, gm_n145);
	or (gm_n1101, gm_n143, in_16, gm_n63, gm_n1100, gm_n237);
	nor (gm_n1102, gm_n89, gm_n82, in_20, gm_n1101, gm_n522);
	nand (gm_n1103, gm_n629, gm_n84, gm_n83, gm_n1102);
	nand (gm_n1104, gm_n1103, gm_n1099, gm_n1095);
	nor (gm_n1105, gm_n1080, gm_n1026, gm_n1022, gm_n1104, gm_n1092);
	and (gm_n1106, gm_n256, gm_n446, gm_n63, gm_n418);
	nand (gm_n1107, gm_n77, in_23, gm_n58, gm_n1106, gm_n455);
	nor (gm_n1108, gm_n612, gm_n55, gm_n54, gm_n1107, gm_n977);
	nor (gm_n1109, gm_n725, in_15, in_11, gm_n503, gm_n669);
	nand (gm_n1110, gm_n74, in_23, in_19, gm_n1109, gm_n173);
	nor (gm_n1111, gm_n57, gm_n55, in_27, gm_n1110, gm_n458);
	not (gm_n1112, gm_n134);
	nor (gm_n1113, gm_n312, gm_n62, gm_n61, gm_n664, gm_n363);
	nand (gm_n1114, gm_n174, in_23, in_19, gm_n1113, gm_n358);
	nor (gm_n1115, gm_n1112, gm_n55, gm_n54, gm_n1114, gm_n838);
	nor (gm_n1116, gm_n1115, gm_n1111, gm_n1108);
	nand (gm_n1117, gm_n515, gm_n311, gm_n124);
	nor (gm_n1118, gm_n188, in_16, gm_n63, gm_n1117, gm_n282);
	nand (gm_n1119, gm_n217, gm_n82, in_20, gm_n1118, gm_n521);
	nor (gm_n1120, gm_n214, gm_n140, gm_n83, gm_n1119);
	nand (gm_n1121, gm_n310, gm_n126, in_11, gm_n502, gm_n426);
	nor (gm_n1122, gm_n131, gm_n58, gm_n62, gm_n1121, gm_n360);
	nand (gm_n1123, gm_n390, gm_n54, gm_n158, gm_n1122, gm_n391);
	nor (gm_n1124, gm_n1123, in_31);
	nor (gm_n1125, in_20, gm_n58, gm_n106);
	nand (gm_n1126, gm_n127, gm_n198, gm_n124, gm_n402);
	nand (gm_n1127, in_12, gm_n61, gm_n66);
	nor (gm_n1128, gm_n534, gm_n105, gm_n175, gm_n1127, gm_n1126);
	nand (gm_n1129, gm_n539, gm_n133, gm_n86, gm_n1128, gm_n1125);
	nor (gm_n1130, in_31, gm_n100, in_29, gm_n1129, gm_n1050);
	nor (gm_n1131, gm_n1130, gm_n1124, gm_n1120);
	nand (gm_n1132, gm_n1105, gm_n1018, gm_n1014, gm_n1131, gm_n1116);
	and (gm_n1133, gm_n731, gm_n189);
	nand (gm_n1134, gm_n126, in_15, in_11, gm_n1133, gm_n931);
	nor (gm_n1135, gm_n431, in_23, in_19, gm_n1134, gm_n393);
	nand (gm_n1136, gm_n308, gm_n55, in_27, gm_n1135, gm_n657);
	nor (gm_n1137, in_2, in_1, gm_n94, in_4, gm_n68);
	nand (gm_n1138, gm_n189, in_12, gm_n124, gm_n1137, gm_n340);
	nor (gm_n1139, gm_n1138, gm_n236);
	and (gm_n1140, gm_n296, gm_n158, gm_n58, gm_n1139, gm_n302);
	nand (gm_n1141, gm_n60, in_31, gm_n54, gm_n1140, gm_n438);
	and (gm_n1142, gm_n515, gm_n219, in_8);
	nand (gm_n1143, gm_n91, gm_n73, gm_n63, gm_n1142, gm_n110);
	nor (gm_n1144, gm_n566, gm_n82, gm_n76, gm_n1143, gm_n463);
	nand (gm_n1145, gm_n139, gm_n81, in_28, gm_n1144);
	nand (gm_n1146, gm_n1145, gm_n1141, gm_n1136);
	nand (gm_n1147, gm_n207, in_16, gm_n63, gm_n913, gm_n228);
	nor (gm_n1148, gm_n197, in_24, in_20, gm_n1147, gm_n104);
	nand (gm_n1149, gm_n339, gm_n101, gm_n83, gm_n1148);
	nor (gm_n1150, gm_n271, gm_n971, in_8);
	nand (gm_n1151, gm_n446, gm_n73, gm_n63, gm_n1150, gm_n242);
	nor (gm_n1152, gm_n187, gm_n82, in_20, gm_n1151, gm_n206);
	nand (gm_n1153, gm_n215, gm_n137, in_28, gm_n1152);
	nor (gm_n1154, gm_n447, gm_n63, in_8, gm_n571, gm_n237);
	nand (gm_n1155, gm_n107, in_20, in_16, gm_n1154, gm_n176);
	nor (gm_n1156, gm_n630, gm_n83, in_24, gm_n1155, gm_n368);
	nand (gm_n1157, gm_n1156, gm_n101);
	nand (gm_n1158, gm_n1157, gm_n1153, gm_n1149);
	nor (gm_n1159, gm_n1132, gm_n1010, gm_n1007, gm_n1158, gm_n1146);
	nand (gm_n1160, gm_n228, gm_n63, gm_n124, gm_n402, gm_n310);
	nor (gm_n1161, gm_n249, gm_n76, in_16, gm_n1160, gm_n476);
	nand (gm_n1162, gm_n215, in_28, gm_n82, gm_n1161, gm_n227);
	nor (gm_n1163, gm_n1162, gm_n479);
	nand (gm_n1164, gm_n453, gm_n218);
	nor (gm_n1165, gm_n553, in_12, in_8, gm_n1164, gm_n352);
	nand (gm_n1166, gm_n235, gm_n76, gm_n73, gm_n1165, gm_n255);
	nor (gm_n1167, gm_n195, gm_n83, in_24, gm_n1166, gm_n262);
	or (gm_n1168, gm_n151, in_6, in_5, gm_n469, in_8);
	nor (gm_n1169, gm_n374, in_16, in_12, gm_n1168, gm_n282);
	nand (gm_n1170, gm_n205, in_24, in_20, gm_n1169, gm_n521);
	nor (gm_n1171, gm_n248, gm_n234, in_28, gm_n1170);
	nor (gm_n1172, gm_n1171, gm_n1167, gm_n1163);
	nor (gm_n1173, gm_n383, gm_n229, gm_n124);
	and (gm_n1174, gm_n200, gm_n73, in_12, gm_n1173, gm_n153);
	nand (gm_n1175, gm_n90, gm_n82, gm_n76, gm_n1174, gm_n205);
	nor (gm_n1176, gm_n195, gm_n224, gm_n83, gm_n1175);
	nor (gm_n1177, gm_n152, gm_n63, gm_n124, gm_n352, gm_n95);
	nor (gm_n1178, gm_n73, in_15, gm_n64);
	and (gm_n1179, gm_n1177, gm_n105, in_13, gm_n1178, gm_n1125);
	nor (gm_n1180, in_24, gm_n158, in_22);
	nand (gm_n1181, gm_n735, gm_n133, gm_n86, gm_n1180, gm_n1179);
	nor (gm_n1182, gm_n55, gm_n100, gm_n80, gm_n1181);
	nor (gm_n1183, gm_n188, in_16, gm_n63, gm_n842, gm_n288);
	nand (gm_n1184, gm_n141, in_24, in_20, gm_n1183, gm_n255);
	nor (gm_n1185, gm_n774, gm_n214, in_28, gm_n1184);
	nor (gm_n1186, gm_n1185, gm_n1182, gm_n1176);
	nand (gm_n1187, gm_n1159, gm_n1003, gm_n999, gm_n1186, gm_n1172);
	or (gm_n1188, gm_n599, in_16, gm_n63, gm_n266, gm_n177);
	nor (gm_n1189, gm_n187, gm_n82, in_20, gm_n1188, gm_n206);
	nand (gm_n1190, gm_n466, gm_n196, in_28, gm_n1189);
	nor (gm_n1191, gm_n92, gm_n63, in_8, gm_n571, gm_n345);
	nand (gm_n1192, gm_n141, gm_n76, in_16, gm_n1191, gm_n150);
	nor (gm_n1193, gm_n85, in_28, in_24, gm_n1192, gm_n206);
	nand (gm_n1194, gm_n1193, gm_n137);
	and (gm_n1195, gm_n620, gm_n144);
	nand (gm_n1196, gm_n300, gm_n62, in_11, gm_n1195, gm_n426);
	nor (gm_n1197, gm_n796, gm_n158, in_19, gm_n1196, gm_n514);
	nand (gm_n1198, gm_n60, gm_n55, in_27, gm_n1197, gm_n511);
	nand (gm_n1199, gm_n1198, gm_n1194, gm_n1190);
	not (gm_n1200, gm_n305);
	nand (gm_n1201, gm_n620, gm_n264);
	nor (gm_n1202, gm_n363, gm_n62, in_11, gm_n1201, gm_n619);
	nand (gm_n1203, gm_n174, gm_n158, gm_n58, gm_n1202, gm_n316);
	nor (gm_n1204, gm_n1200, in_31, in_27, gm_n1203, gm_n612);
	nor (out_3, gm_n1199, gm_n1187, gm_n994, gm_n1204);
	and (gm_n1206, gm_n207, in_20, gm_n73, gm_n1154, gm_n477);
	nand (gm_n1207, gm_n103, gm_n83, gm_n82, gm_n1206, gm_n466);
	nor (gm_n1208, gm_n1207, gm_n185);
	nand (gm_n1209, gm_n402, gm_n264);
	or (gm_n1210, gm_n249, in_12, gm_n124, gm_n1209, gm_n237);
	nor (gm_n1211, gm_n801, in_20, in_16, gm_n1210, gm_n522);
	nand (gm_n1212, gm_n186, in_28, in_24, gm_n1211, gm_n225);
	and (gm_n1213, gm_n167, in_12, in_8, gm_n515, gm_n243);
	nand (gm_n1214, gm_n142, gm_n76, in_16, gm_n1213, gm_n270);
	nor (gm_n1215, gm_n85, gm_n83, gm_n82, gm_n1214, gm_n89);
	nand (gm_n1216, gm_n1215, gm_n196);
	nand (gm_n1217, gm_n151, in_6, in_5, gm_n361, in_8);
	nor (gm_n1218, gm_n249, in_16, gm_n63, gm_n1217, gm_n237);
	nand (gm_n1219, gm_n90, gm_n82, gm_n76, gm_n1218, gm_n217);
	nor (gm_n1220, gm_n368, gm_n214, in_28, gm_n1219);
	nand (gm_n1221, gm_n594, gm_n515);
	nor (gm_n1222, gm_n322, gm_n62, in_11, gm_n1221, gm_n425);
	nand (gm_n1223, gm_n174, in_23, in_19, gm_n1222, gm_n296);
	nor (gm_n1224, gm_n357, gm_n55, in_27, gm_n1223, gm_n583);
	not (gm_n1225, gm_n77);
	not (gm_n1226, gm_n991);
	nand (gm_n1227, gm_n72, in_15, in_11, gm_n1226, gm_n392);
	nor (gm_n1228, gm_n1225, in_23, gm_n58, gm_n1227, gm_n1200);
	nand (gm_n1229, gm_n337, gm_n55, in_27, gm_n1228);
	nand (gm_n1230, gm_n243, gm_n189, in_8);
	or (gm_n1231, gm_n249, in_16, in_12, gm_n1230, gm_n154);
	nor (gm_n1232, gm_n89, gm_n82, gm_n76, gm_n1231, gm_n187);
	nand (gm_n1233, gm_n215, gm_n81, gm_n83, gm_n1232);
	or (gm_n1234, gm_n345, gm_n114, in_8);
	nor (gm_n1235, gm_n249, gm_n73, gm_n63, gm_n1234, gm_n111);
	nand (gm_n1236, gm_n205, in_24, in_20, gm_n1235, gm_n235);
	nor (gm_n1237, gm_n684, gm_n368, gm_n83, gm_n1236);
	nor (gm_n1238, gm_n92, gm_n63, gm_n124, gm_n965, gm_n553);
	nand (gm_n1239, gm_n164, in_20, in_16, gm_n1238, gm_n227);
	nor (gm_n1240, gm_n138, in_28, in_24, gm_n1239, gm_n262);
	nand (gm_n1241, gm_n110, in_16, in_12, gm_n1011, gm_n207);
	nor (gm_n1242, gm_n566, gm_n82, in_20, gm_n1241, gm_n522);
	nand (gm_n1243, gm_n225, gm_n139, gm_n83, gm_n1242);
	nand (gm_n1244, in_5, in_4, gm_n68, gm_n145, gm_n115);
	nor (gm_n1245, gm_n1244, in_8, in_7);
	nand (gm_n1246, gm_n166, in_16, in_12, gm_n1245, gm_n167);
	nor (gm_n1247, gm_n197, in_24, gm_n76, gm_n1246, gm_n206);
	nand (gm_n1248, gm_n466, gm_n196, gm_n83, gm_n1247);
	nor (gm_n1249, gm_n363, gm_n62, in_11, gm_n726, gm_n664);
	nand (gm_n1250, gm_n358, in_23, gm_n58, gm_n1249, gm_n359);
	nor (gm_n1251, gm_n422, in_31, gm_n54, gm_n1250, gm_n612);
	nand (gm_n1252, gm_n453, gm_n264);
	nor (gm_n1253, gm_n432, gm_n62, gm_n61, gm_n1252, gm_n664);
	nand (gm_n1254, gm_n130, in_23, in_19, gm_n1253, gm_n455);
	nor (gm_n1255, gm_n423, in_31, gm_n54, gm_n1254, gm_n977);
	nor (gm_n1256, gm_n553, in_12, in_8, gm_n554, gm_n352);
	nand (gm_n1257, gm_n192, gm_n76, in_16, gm_n1256, gm_n235);
	nor (gm_n1258, gm_n138, in_28, in_24, gm_n1257, gm_n368);
	or (gm_n1259, gm_n151, gm_n115, gm_n70, gm_n168);
	nor (gm_n1260, gm_n664, gm_n62, gm_n61, gm_n1259, gm_n991);
	nand (gm_n1261, gm_n173, gm_n158, in_19, gm_n1260, gm_n455);
	nor (gm_n1262, gm_n357, in_31, in_27, gm_n1261, gm_n583);
	or (gm_n1263, gm_n971, gm_n114, gm_n124);
	nor (gm_n1264, gm_n374, in_16, in_12, gm_n1263, gm_n352);
	nand (gm_n1265, gm_n103, in_24, in_20, gm_n1264, gm_n107);
	nor (gm_n1266, gm_n262, gm_n214, in_28, gm_n1265);
	nor (gm_n1267, gm_n1258, gm_n1255, gm_n1251, gm_n1266, gm_n1262);
	nand (gm_n1268, gm_n243, gm_n71);
	nor (gm_n1269, gm_n669, in_15, in_11, gm_n1268, gm_n670);
	nand (gm_n1270, gm_n174, in_23, in_19, gm_n1269, gm_n316);
	nor (gm_n1271, gm_n583, gm_n55, gm_n54, gm_n1270, gm_n838);
	nand (gm_n1272, gm_n115, gm_n70, gm_n113, gm_n543, gm_n151);
	nor (gm_n1273, gm_n125, in_15, gm_n61, gm_n1272, gm_n314);
	nand (gm_n1274, gm_n77, gm_n158, in_19, gm_n1273, gm_n359);
	nor (gm_n1275, gm_n618, gm_n55, in_27, gm_n1274, gm_n977);
	nand (gm_n1276, gm_n515, gm_n128);
	nor (gm_n1277, gm_n177, gm_n63, gm_n124, gm_n1276, gm_n237);
	nand (gm_n1278, gm_n174, in_23, in_19, gm_n1277, gm_n358);
	nor (gm_n1279, gm_n1112, gm_n55, gm_n54, gm_n1278, gm_n612);
	nor (gm_n1280, gm_n1279, gm_n1275, gm_n1271);
	and (gm_n1281, gm_n200, in_16, gm_n63, gm_n887, gm_n256);
	nand (gm_n1282, gm_n107, in_24, in_20, gm_n1281, gm_n205);
	nor (gm_n1283, gm_n138, gm_n224, gm_n83, gm_n1282);
	nor (gm_n1284, gm_n143, gm_n73, in_12, gm_n905, gm_n237);
	nand (gm_n1285, gm_n90, in_24, gm_n76, gm_n1284, gm_n192);
	nor (gm_n1286, gm_n479, gm_n248, in_28, gm_n1285);
	nand (gm_n1287, in_7, gm_n115, gm_n70, gm_n361, gm_n124);
	nor (gm_n1288, gm_n236, gm_n73, gm_n63, gm_n1287, gm_n599);
	nand (gm_n1289, gm_n205, in_24, in_20, gm_n1288, gm_n477);
	nor (gm_n1290, gm_n224, gm_n234, in_28, gm_n1289);
	nor (gm_n1291, gm_n1290, gm_n1286, gm_n1283);
	nand (gm_n1292, gm_n1267, gm_n1248, gm_n1243, gm_n1291, gm_n1280);
	nand (gm_n1293, gm_n199, in_16, gm_n63, gm_n272, gm_n150);
	nor (gm_n1294, gm_n104, in_24, in_20, gm_n1293, gm_n187);
	nand (gm_n1295, gm_n466, gm_n225, in_28, gm_n1294);
	nand (gm_n1296, gm_n775, gm_n264, in_8);
	or (gm_n1297, gm_n143, in_16, gm_n63, gm_n1296, gm_n282);
	nor (gm_n1298, gm_n89, gm_n82, in_20, gm_n1297, gm_n412);
	nand (gm_n1299, gm_n367, gm_n196, gm_n83, gm_n1298);
	nor (gm_n1300, gm_n116, gm_n63, in_8, gm_n288, gm_n972);
	nand (gm_n1301, gm_n141, gm_n76, gm_n73, gm_n1300, gm_n150);
	nor (gm_n1302, gm_n262, in_28, in_24, gm_n1301, gm_n630);
	nand (gm_n1303, gm_n1302, gm_n629);
	nand (gm_n1304, gm_n1303, gm_n1299, gm_n1295);
	nand (gm_n1305, gm_n91, in_16, gm_n63, gm_n516, gm_n199);
	nor (gm_n1306, gm_n104, in_24, gm_n76, gm_n1305, gm_n108);
	nand (gm_n1307, gm_n137, gm_n84, in_28, gm_n1306);
	and (gm_n1308, gm_n189, gm_n63, in_8, gm_n588, gm_n167);
	nand (gm_n1309, gm_n207, gm_n76, gm_n73, gm_n1308, gm_n235);
	nor (gm_n1310, gm_n520, gm_n83, gm_n82, gm_n1309, gm_n368);
	nand (gm_n1311, gm_n1310, gm_n225);
	and (gm_n1312, gm_n453, gm_n144);
	nand (gm_n1313, gm_n426, gm_n62, gm_n61, gm_n1312, gm_n730);
	nor (gm_n1314, gm_n122, in_23, gm_n58, gm_n1313, gm_n131);
	nand (gm_n1315, gm_n309, in_31, gm_n54, gm_n1314, gm_n511);
	nand (gm_n1316, gm_n1315, gm_n1311, gm_n1307);
	nor (gm_n1317, gm_n1292, gm_n1240, gm_n1237, gm_n1316, gm_n1304);
	nand (gm_n1318, gm_n218, gm_n69, in_8);
	nor (gm_n1319, gm_n92, in_16, in_12, gm_n1318, gm_n143);
	nand (gm_n1320, gm_n263, in_24, gm_n76, gm_n1319, gm_n521);
	nor (gm_n1321, gm_n248, gm_n234, in_28, gm_n1320);
	nand (gm_n1322, gm_n594, gm_n189);
	nor (gm_n1323, gm_n314, gm_n62, in_11, gm_n1322, gm_n619);
	nand (gm_n1324, gm_n74, in_23, in_19, gm_n1323, gm_n77);
	nor (gm_n1325, gm_n57, gm_n55, gm_n54, gm_n1324, gm_n458);
	or (gm_n1326, gm_n152, gm_n63, gm_n124, gm_n288, gm_n95);
	nor (gm_n1327, gm_n197, gm_n76, in_16, gm_n1326, gm_n236);
	nand (gm_n1328, gm_n215, in_28, gm_n82, gm_n1327, gm_n255);
	nor (gm_n1329, gm_n1328, gm_n234);
	nor (gm_n1330, gm_n1329, gm_n1325, gm_n1321);
	nor (gm_n1331, in_7, gm_n115, in_5, gm_n469, in_8);
	and (gm_n1332, gm_n153, in_16, in_12, gm_n1331, gm_n207);
	nand (gm_n1333, gm_n255, gm_n82, in_20, gm_n1332, gm_n270);
	nor (gm_n1334, gm_n138, gm_n85, in_28, gm_n1333);
	and (gm_n1335, gm_n207, in_16, in_12, gm_n572, gm_n256);
	nand (gm_n1336, gm_n192, in_24, gm_n76, gm_n1335, gm_n477);
	nor (gm_n1337, gm_n684, gm_n224, in_28, gm_n1336);
	nor (gm_n1338, gm_n321, in_15, gm_n61, gm_n425, gm_n433);
	nand (gm_n1339, gm_n121, gm_n158, gm_n58, gm_n1338, gm_n358);
	nor (gm_n1340, gm_n357, in_31, gm_n54, gm_n1339, gm_n977);
	nor (gm_n1341, gm_n1340, gm_n1337, gm_n1334);
	nand (gm_n1342, gm_n1317, gm_n1233, gm_n1229, gm_n1341, gm_n1330);
	or (gm_n1343, gm_n109, in_16, gm_n63, gm_n905, gm_n111);
	nor (gm_n1344, gm_n197, gm_n82, gm_n76, gm_n1343, gm_n801);
	nand (gm_n1345, gm_n215, gm_n101, gm_n83, gm_n1344);
	nor (gm_n1346, gm_n447, gm_n63, gm_n124, gm_n229, gm_n599);
	nand (gm_n1347, gm_n90, in_20, in_16, gm_n1346, gm_n91);
	nor (gm_n1348, gm_n224, in_28, in_24, gm_n1347, gm_n801);
	nand (gm_n1349, gm_n1348, gm_n101);
	and (gm_n1350, gm_n502, gm_n264, gm_n124);
	nand (gm_n1351, gm_n153, gm_n73, in_12, gm_n1350, gm_n207);
	nor (gm_n1352, gm_n520, in_24, gm_n76, gm_n1351, gm_n476);
	nand (gm_n1353, gm_n629, gm_n367, gm_n83, gm_n1352);
	nand (gm_n1354, gm_n1353, gm_n1349, gm_n1345);
	and (gm_n1355, gm_n264, gm_n243, gm_n124);
	nand (gm_n1356, gm_n176, in_16, gm_n63, gm_n1355, gm_n256);
	nor (gm_n1357, gm_n187, in_24, gm_n76, gm_n1356, gm_n520);
	nand (gm_n1358, gm_n102, gm_n81, gm_n83, gm_n1357);
	nand (gm_n1359, gm_n703, gm_n264, gm_n124);
	or (gm_n1360, gm_n111, in_16, gm_n63, gm_n1359, gm_n236);
	nor (gm_n1361, gm_n206, gm_n82, gm_n76, gm_n1360, gm_n463);
	nand (gm_n1362, gm_n139, gm_n81, gm_n83, gm_n1361);
	nor (gm_n1363, gm_n151, in_6, gm_n70, gm_n469, gm_n124);
	nand (gm_n1364, gm_n150, gm_n73, in_12, gm_n1363, gm_n340);
	nor (gm_n1365, gm_n104, gm_n82, gm_n76, gm_n1364, gm_n522);
	nand (gm_n1366, gm_n339, gm_n101, in_28, gm_n1365);
	nand (gm_n1367, gm_n1366, gm_n1362, gm_n1358);
	nor (gm_n1368, gm_n1342, gm_n1224, gm_n1220, gm_n1367, gm_n1354);
	nor (gm_n1369, gm_n188, in_12, gm_n124, gm_n288, gm_n284);
	nand (gm_n1370, gm_n141, gm_n76, in_16, gm_n1369, gm_n205);
	nor (gm_n1371, gm_n248, in_28, gm_n82, gm_n1370, gm_n226);
	nor (gm_n1372, gm_n177, in_16, gm_n63, gm_n654, gm_n282);
	nand (gm_n1373, gm_n192, in_24, in_20, gm_n1372, gm_n477);
	nor (gm_n1374, gm_n479, gm_n368, gm_n83, gm_n1373);
	nor (gm_n1375, gm_n553, gm_n73, gm_n63, gm_n1100, gm_n282);
	nand (gm_n1376, gm_n90, in_24, gm_n76, gm_n1375, gm_n217);
	nor (gm_n1377, gm_n248, gm_n234, gm_n83, gm_n1376);
	nor (gm_n1378, gm_n1377, gm_n1374, gm_n1371);
	nand (gm_n1379, gm_n69, in_12, in_8, gm_n264, gm_n199);
	nor (gm_n1380, gm_n177, gm_n76, gm_n73, gm_n1379, gm_n412);
	nand (gm_n1381, gm_n186, in_28, in_24, gm_n1380, gm_n263);
	nor (gm_n1382, gm_n1381, gm_n234);
	or (gm_n1383, gm_n469, gm_n383, in_8);
	nor (gm_n1384, gm_n177, in_16, gm_n63, gm_n1383, gm_n282);
	nand (gm_n1385, gm_n263, gm_n82, in_20, gm_n1384, gm_n477);
	nor (gm_n1386, gm_n214, gm_n248, gm_n83, gm_n1385);
	nand (gm_n1387, gm_n283, gm_n127, gm_n124);
	nor (gm_n1388, gm_n249, gm_n73, in_12, gm_n1387, gm_n599);
	nand (gm_n1389, gm_n164, in_24, gm_n76, gm_n1388, gm_n227);
	nor (gm_n1390, gm_n684, gm_n368, gm_n83, gm_n1389);
	nor (gm_n1391, gm_n1390, gm_n1386, gm_n1382);
	nand (gm_n1392, gm_n1368, gm_n1216, gm_n1212, gm_n1391, gm_n1378);
	and (gm_n1393, gm_n123, gm_n71, in_11, gm_n502, gm_n394);
	nand (gm_n1394, gm_n302, gm_n58, gm_n62, gm_n1393, gm_n334);
	nor (gm_n1395, gm_n423, in_27, in_23, gm_n1394, gm_n977);
	nand (gm_n1396, gm_n1395, in_31);
	nand (gm_n1397, gm_n930, gm_n62, in_11, gm_n792, gm_n426);
	nor (gm_n1398, gm_n796, in_23, gm_n58, gm_n1397, gm_n431);
	nand (gm_n1399, gm_n309, in_31, gm_n54, gm_n1398, gm_n337);
	and (gm_n1400, gm_n311, gm_n144);
	nand (gm_n1401, gm_n698, in_15, in_11, gm_n1400, gm_n424);
	nor (gm_n1402, gm_n122, gm_n158, in_19, gm_n1401, gm_n452);
	nand (gm_n1403, gm_n308, in_31, in_27, gm_n1402, gm_n657);
	nand (gm_n1404, gm_n1403, gm_n1399, gm_n1396);
	nand (gm_n1405, gm_n265, gm_n218, gm_n124);
	nor (gm_n1406, gm_n143, gm_n73, in_12, gm_n1405, gm_n154);
	nand (gm_n1407, gm_n164, in_24, gm_n76, gm_n1406, gm_n227);
	nor (gm_n1408, gm_n368, gm_n185, in_28, gm_n1407);
	nor (out_4, gm_n1404, gm_n1392, gm_n1208, gm_n1408);
	nand (gm_n1410, gm_n167, gm_n63, gm_n124, gm_n402, gm_n515);
	nor (gm_n1411, gm_n108, in_20, in_16, gm_n1410, gm_n177);
	nand (gm_n1412, gm_n263, gm_n83, gm_n82, gm_n1411, gm_n367);
	nor (gm_n1413, gm_n1412, gm_n138);
	nand (gm_n1414, gm_n107, in_20, gm_n73, gm_n957, gm_n142);
	nor (gm_n1415, gm_n85, gm_n83, gm_n82, gm_n1414, gm_n206);
	nand (gm_n1416, gm_n1415, gm_n629);
	nor (gm_n1417, gm_n152, in_12, in_8, gm_n599, gm_n95);
	nand (gm_n1418, gm_n141, in_20, gm_n73, gm_n1417, gm_n176);
	nor (gm_n1419, gm_n224, gm_n83, in_24, gm_n1418, gm_n206);
	nand (gm_n1420, gm_n1419, gm_n496);
	nand (gm_n1421, gm_n110, in_12, gm_n124, gm_n243, gm_n189);
	nor (gm_n1422, gm_n236, gm_n76, in_16, gm_n1421, gm_n522);
	nand (gm_n1423, gm_n102, in_28, in_24, gm_n1422, gm_n227);
	nor (gm_n1424, gm_n1423, gm_n138);
	nand (gm_n1425, gm_n218, in_12, in_8, gm_n703, gm_n167);
	nor (gm_n1426, gm_n249, in_20, gm_n73, gm_n1425, gm_n476);
	nand (gm_n1427, gm_n103, gm_n83, in_24, gm_n1426, gm_n215);
	nor (gm_n1428, gm_n1427, gm_n195);
	or (gm_n1429, gm_n177, in_16, in_12, gm_n1063, gm_n237);
	nor (gm_n1430, gm_n104, gm_n82, gm_n76, gm_n1429, gm_n412);
	nand (gm_n1431, gm_n186, gm_n137, gm_n83, gm_n1430);
	and (gm_n1432, gm_n144, in_12, in_8, gm_n588, gm_n242);
	nand (gm_n1433, gm_n107, in_20, in_16, gm_n1432, gm_n142);
	nor (gm_n1434, gm_n216, in_28, in_24, gm_n1433, gm_n630);
	nand (gm_n1435, gm_n1434, gm_n496);
	nor (gm_n1436, gm_n553, gm_n73, gm_n63, gm_n1383, gm_n288);
	nand (gm_n1437, gm_n217, gm_n82, gm_n76, gm_n1436, gm_n270);
	nor (gm_n1438, gm_n195, gm_n248, in_28, gm_n1437);
	nand (gm_n1439, gm_n69, in_12, gm_n124, gm_n515, gm_n199);
	nor (gm_n1440, gm_n249, in_20, gm_n73, gm_n1439, gm_n108);
	nand (gm_n1441, gm_n84, gm_n83, in_24, gm_n1440, gm_n217);
	nor (gm_n1442, gm_n1441, gm_n195);
	nand (gm_n1443, gm_n1042, in_15, gm_n61, gm_n1226, gm_n948);
	nor (gm_n1444, gm_n1112, in_23, gm_n58, gm_n1443, gm_n431);
	nand (gm_n1445, gm_n306, gm_n55, gm_n54, gm_n1444);
	nand (gm_n1446, gm_n446, in_16, in_12, gm_n346, gm_n228);
	nor (gm_n1447, gm_n89, gm_n82, gm_n76, gm_n1446, gm_n108);
	nand (gm_n1448, gm_n466, gm_n196, in_28, gm_n1447);
	nor (gm_n1449, gm_n143, in_16, gm_n63, gm_n1063, gm_n288);
	nand (gm_n1450, gm_n255, gm_n82, gm_n76, gm_n1449, gm_n521);
	nor (gm_n1451, gm_n216, gm_n214, gm_n83, gm_n1450);
	and (gm_n1452, gm_n153, gm_n142, in_12, gm_n1042, gm_n589);
	nand (gm_n1453, gm_n296, gm_n158, in_19, gm_n1452, gm_n657);
	nor (gm_n1454, gm_n437, in_31, in_27, gm_n1453);
	nor (gm_n1455, gm_n284, in_15, in_11, gm_n619, gm_n314);
	nand (gm_n1456, gm_n173, gm_n158, in_19, gm_n1455, gm_n392);
	nor (gm_n1457, gm_n618, in_31, gm_n54, gm_n1456, gm_n583);
	and (gm_n1458, gm_n110, in_16, gm_n63, gm_n883, gm_n207);
	nand (gm_n1459, gm_n88, gm_n82, in_20, gm_n1458, gm_n164);
	nor (gm_n1460, gm_n214, gm_n140, gm_n83, gm_n1459);
	nor (gm_n1461, gm_n249, gm_n73, gm_n63, gm_n1068, gm_n352);
	nand (gm_n1462, gm_n192, gm_n82, gm_n76, gm_n1461, gm_n521);
	nor (gm_n1463, gm_n262, gm_n138, in_28, gm_n1462);
	nor (gm_n1464, gm_n1457, gm_n1454, gm_n1451, gm_n1463, gm_n1460);
	nand (gm_n1465, gm_n310, gm_n340, gm_n124, gm_n731, gm_n426);
	nor (gm_n1466, gm_n297, in_19, gm_n62, gm_n1465, gm_n613);
	nand (gm_n1467, gm_n60, gm_n54, in_23, gm_n1466, gm_n674);
	nor (gm_n1468, gm_n1467, in_31);
	nor (gm_n1469, gm_n122, gm_n62, gm_n61, gm_n362, gm_n669);
	nand (gm_n1470, gm_n77, in_23, in_19, gm_n1469, gm_n391);
	nor (gm_n1471, gm_n57, gm_n55, in_27, gm_n1470);
	nor (gm_n1472, gm_n109, in_16, gm_n63, gm_n1234, gm_n154);
	nand (gm_n1473, gm_n227, gm_n82, in_20, gm_n1472, gm_n477);
	nor (gm_n1474, gm_n479, gm_n216, in_28, gm_n1473);
	nor (gm_n1475, gm_n1474, gm_n1471, gm_n1468);
	nor (gm_n1476, gm_n92, gm_n63, in_8, gm_n1276, gm_n177);
	nand (gm_n1477, gm_n205, gm_n76, gm_n73, gm_n1476, gm_n270);
	nor (gm_n1478, gm_n140, in_28, in_24, gm_n1477, gm_n479);
	nand (gm_n1479, gm_n219, gm_n127);
	nor (gm_n1480, gm_n322, gm_n62, in_11, gm_n1479, gm_n363);
	nand (gm_n1481, gm_n173, gm_n158, in_19, gm_n1480, gm_n1042);
	nor (gm_n1482, gm_n183, in_31, in_27, gm_n1481, gm_n437);
	nor (gm_n1483, gm_n143, in_12, gm_n124, gm_n1209, gm_n154);
	nand (gm_n1484, gm_n217, in_20, gm_n73, gm_n1483, gm_n270);
	nor (gm_n1485, gm_n224, gm_n83, in_24, gm_n1484, gm_n479);
	nor (gm_n1486, gm_n1485, gm_n1482, gm_n1478);
	nand (gm_n1487, gm_n1464, gm_n1448, gm_n1445, gm_n1486, gm_n1475);
	nand (gm_n1488, gm_n313, gm_n153, in_15, gm_n1142, gm_n455);
	nor (gm_n1489, gm_n422, gm_n158, gm_n58, gm_n1488, gm_n317);
	nand (gm_n1490, gm_n390, gm_n55, in_27, gm_n1489);
	and (gm_n1491, gm_n264, gm_n69, gm_n124);
	nand (gm_n1492, gm_n199, in_16, in_12, gm_n1491, gm_n142);
	nor (gm_n1493, gm_n197, gm_n82, gm_n76, gm_n1492, gm_n411);
	nand (gm_n1494, gm_n466, gm_n225, gm_n83, gm_n1493);
	nand (gm_n1495, gm_n176, in_16, in_12, gm_n470, gm_n242);
	nor (gm_n1496, gm_n108, gm_n82, gm_n76, gm_n1495, gm_n630);
	nand (gm_n1497, gm_n102, gm_n81, in_28, gm_n1496);
	nand (gm_n1498, gm_n1497, gm_n1494, gm_n1490);
	and (gm_n1499, gm_n453, gm_n144, gm_n124);
	nand (gm_n1500, gm_n110, in_16, in_12, gm_n1499, gm_n150);
	nor (gm_n1501, gm_n520, in_24, in_20, gm_n1500, gm_n412);
	nand (gm_n1502, gm_n339, gm_n213, gm_n83, gm_n1501);
	or (gm_n1503, gm_n146, in_12, in_8, gm_n237, gm_n553);
	nor (gm_n1504, gm_n520, in_20, gm_n73, gm_n1503, gm_n476);
	nand (gm_n1505, gm_n137, in_28, gm_n82, gm_n1504, gm_n367);
	and (gm_n1506, gm_n310, gm_n243);
	nand (gm_n1507, gm_n167, in_12, in_8, gm_n1506, gm_n207);
	nor (gm_n1508, gm_n104, in_20, in_16, gm_n1507, gm_n522);
	nand (gm_n1509, gm_n101, in_28, gm_n82, gm_n1508, gm_n466);
	nand (gm_n1510, gm_n1509, gm_n1505, gm_n1502);
	nor (gm_n1511, gm_n1487, gm_n1442, gm_n1438, gm_n1510, gm_n1498);
	nand (gm_n1512, gm_n731, gm_n515);
	nor (gm_n1513, gm_n619, gm_n62, in_11, gm_n1512, gm_n623);
	nand (gm_n1514, gm_n77, gm_n158, gm_n58, gm_n1513, gm_n455);
	nor (gm_n1515, gm_n357, in_31, gm_n54, gm_n1514, gm_n422);
	nor (gm_n1516, gm_n108, in_20, gm_n73, gm_n818, gm_n553);
	nand (gm_n1517, gm_n84, in_28, in_24, gm_n1516, gm_n217);
	nor (gm_n1518, gm_n1517, gm_n195);
	nand (gm_n1519, gm_n775, gm_n218, in_8);
	nor (gm_n1520, gm_n154, gm_n73, gm_n63, gm_n1519, gm_n177);
	nand (gm_n1521, gm_n88, gm_n82, gm_n76, gm_n1520, gm_n107);
	nor (gm_n1522, gm_n214, gm_n140, in_28, gm_n1521);
	nor (gm_n1523, gm_n1522, gm_n1518, gm_n1515);
	nor (gm_n1524, gm_n393, in_19, gm_n62, gm_n996, gm_n991);
	nand (gm_n1525, gm_n358, gm_n54, in_23, gm_n1524, gm_n657);
	nor (gm_n1526, gm_n1525, gm_n618, gm_n55);
	nand (gm_n1527, gm_n310, gm_n396);
	nor (gm_n1528, gm_n669, gm_n62, gm_n124, gm_n1527, gm_n288);
	nand (gm_n1529, gm_n173, gm_n158, in_19, gm_n1528, gm_n455);
	nor (gm_n1530, gm_n458, gm_n55, in_27, gm_n1529, gm_n675);
	nand (gm_n1531, gm_n588, gm_n424, gm_n189);
	nor (gm_n1532, gm_n796, in_15, gm_n61, gm_n1531, gm_n669);
	nand (gm_n1533, gm_n130, in_23, gm_n58, gm_n1532, gm_n309);
	nor (gm_n1534, gm_n437, in_31, gm_n54, gm_n1533);
	nor (gm_n1535, gm_n1534, gm_n1530, gm_n1526);
	nand (gm_n1536, gm_n1511, gm_n1435, gm_n1431, gm_n1535, gm_n1523);
	nor (gm_n1537, gm_n151, in_6, in_5, gm_n469);
	nand (gm_n1538, gm_n65, in_15, gm_n61, gm_n1537, gm_n797);
	nor (gm_n1539, gm_n431, gm_n158, in_19, gm_n1538, gm_n360);
	nand (gm_n1540, gm_n657, in_31, in_27, gm_n1539, gm_n674);
	nand (gm_n1541, gm_n124, gm_n113, gm_n68, gm_n145, gm_n218);
	or (gm_n1542, gm_n143, in_16, in_12, gm_n1541, gm_n352);
	nor (gm_n1543, gm_n197, in_24, gm_n76, gm_n1542, gm_n630);
	nand (gm_n1544, gm_n629, gm_n139, gm_n83, gm_n1543);
	and (gm_n1545, gm_n730, gm_n310, gm_n208);
	nand (gm_n1546, gm_n121, gm_n62, gm_n61, gm_n1545, gm_n123);
	nor (gm_n1547, gm_n183, gm_n158, in_19, gm_n1546, gm_n514);
	nand (gm_n1548, gm_n308, gm_n55, gm_n54, gm_n1547);
	nand (gm_n1549, gm_n1548, gm_n1544, gm_n1540);
	or (gm_n1550, gm_n669, in_15, in_11, gm_n584, gm_n670);
	nor (gm_n1551, gm_n331, gm_n158, gm_n58, gm_n1550, gm_n335);
	nand (gm_n1552, gm_n306, gm_n55, gm_n54, gm_n1551, gm_n459);
	and (gm_n1553, gm_n620, gm_n127, in_8);
	nand (gm_n1554, gm_n91, gm_n73, gm_n63, gm_n1553, gm_n228);
	nor (gm_n1555, gm_n566, gm_n82, gm_n76, gm_n1554, gm_n476);
	nand (gm_n1556, gm_n225, gm_n84, gm_n83, gm_n1555);
	not (gm_n1557, gm_n326);
	nor (gm_n1558, gm_n152, gm_n198, gm_n124, gm_n753);
	nand (gm_n1559, gm_n63, gm_n61, gm_n66, gm_n1558, gm_n175);
	nor (gm_n1560, in_20, in_19, in_18);
	not (gm_n1561, gm_n1560);
	or (gm_n1562, gm_n767, gm_n86, gm_n105, gm_n1561, gm_n1559);
	nor (gm_n1563, gm_n1562, gm_n1557, in_25);
	nand (gm_n1564, gm_n55, in_30, gm_n80, gm_n1563, gm_n540);
	nand (gm_n1565, gm_n1564, gm_n1556, gm_n1552);
	nor (gm_n1566, gm_n1536, gm_n1428, gm_n1424, gm_n1565, gm_n1549);
	nor (gm_n1567, gm_n360, gm_n237, in_15, gm_n1046, gm_n363);
	nand (gm_n1568, gm_n130, gm_n158, gm_n58, gm_n1567, gm_n182);
	nor (gm_n1569, gm_n437, in_31, in_27, gm_n1568);
	nand (gm_n1570, gm_n144, gm_n63, gm_n124, gm_n243, gm_n153);
	nor (gm_n1571, gm_n1570, gm_n188, in_16);
	nand (gm_n1572, gm_n227, gm_n82, gm_n76, gm_n1571, gm_n477);
	nor (gm_n1573, gm_n140, gm_n138, in_28, gm_n1572);
	nor (gm_n1574, gm_n271, gm_n93, gm_n124);
	and (gm_n1575, gm_n166, in_16, gm_n63, gm_n1574, gm_n167);
	nand (gm_n1576, gm_n255, in_24, gm_n76, gm_n1575, gm_n270);
	nor (gm_n1577, gm_n226, gm_n140, gm_n83, gm_n1576);
	nor (gm_n1578, gm_n1577, gm_n1573, gm_n1569);
	nor (gm_n1579, gm_n395, in_15, in_11, gm_n1512, gm_n425);
	nand (gm_n1580, gm_n77, gm_n158, gm_n58, gm_n1579, gm_n302);
	nor (gm_n1581, gm_n57, gm_n55, in_27, gm_n1580, gm_n183);
	nor (gm_n1582, gm_n154, in_16, in_12, gm_n1023, gm_n177);
	nand (gm_n1583, gm_n192, in_24, in_20, gm_n1582, gm_n521);
	nor (gm_n1584, gm_n479, gm_n248, gm_n83, gm_n1583);
	nor (gm_n1585, gm_n177, gm_n73, gm_n63, gm_n631, gm_n288);
	nand (gm_n1586, gm_n90, gm_n82, gm_n76, gm_n1585, gm_n255);
	nor (gm_n1587, gm_n774, gm_n195, gm_n83, gm_n1586);
	nor (gm_n1588, gm_n1587, gm_n1584, gm_n1581);
	nand (gm_n1589, gm_n1566, gm_n1420, gm_n1416, gm_n1588, gm_n1578);
	nor (gm_n1590, gm_n178, gm_n152, gm_n124);
	nand (gm_n1591, gm_n110, in_16, in_12, gm_n1590, gm_n446);
	nor (gm_n1592, gm_n630, in_24, in_20, gm_n1591, gm_n522);
	nand (gm_n1593, gm_n139, gm_n137, gm_n83, gm_n1592);
	nand (gm_n1594, gm_n153, gm_n123, gm_n62, gm_n1142, gm_n174);
	nor (gm_n1595, gm_n335, gm_n158, gm_n58, gm_n1594, gm_n583);
	nand (gm_n1596, gm_n390, in_31, gm_n54, gm_n1595);
	and (gm_n1597, gm_n180, gm_n158, gm_n58, gm_n455, gm_n334);
	nand (gm_n1598, gm_n182, in_31, gm_n54, gm_n1597, gm_n511);
	nand (gm_n1599, gm_n1598, gm_n1596, gm_n1593);
	nor (gm_n1600, gm_n143, gm_n73, gm_n63, gm_n1318, gm_n599);
	nand (gm_n1601, gm_n205, in_24, in_20, gm_n1600, gm_n270);
	nor (gm_n1602, gm_n368, gm_n226, in_28, gm_n1601);
	nor (out_5, gm_n1599, gm_n1589, gm_n1413, gm_n1602);
	nor (gm_n1604, gm_n198, gm_n124, in_7);
	and (gm_n1605, in_5, in_4, gm_n68, gm_n145, gm_n115);
	nand (gm_n1606, gm_n636, gm_n1604, gm_n66, gm_n1605);
	nor (gm_n1607, gm_n534, gm_n86, in_17, gm_n1606, gm_n1561);
	nand (gm_n1608, gm_n326, gm_n80, gm_n133, gm_n1607, gm_n735);
	nor (gm_n1609, gm_n1608, gm_n55, gm_n100);
	nand (gm_n1610, gm_n200, in_16, in_12, gm_n1245, gm_n153);
	nor (gm_n1611, gm_n197, in_24, in_20, gm_n1610, gm_n801);
	nand (gm_n1612, gm_n186, gm_n81, in_28, gm_n1611);
	nand (gm_n1613, in_9, gm_n124, in_7);
	nor (gm_n1614, gm_n63, gm_n61, gm_n66, gm_n1613, gm_n1244);
	nand (gm_n1615, gm_n1614, gm_n150);
	nor (gm_n1616, gm_n331, gm_n158, gm_n58, gm_n1615, gm_n335);
	nand (gm_n1617, gm_n309, in_31, gm_n54, gm_n1616, gm_n337);
	or (gm_n1618, gm_n548, gm_n447, gm_n125);
	nor (gm_n1619, gm_n331, gm_n62, in_11, gm_n1618, gm_n623);
	nand (gm_n1620, gm_n173, in_23, in_19, gm_n1619, gm_n459);
	nor (gm_n1621, gm_n423, gm_n55, in_27, gm_n1620);
	or (gm_n1622, gm_n114, gm_n93, in_11, gm_n623, gm_n322);
	nor (gm_n1623, gm_n122, in_19, in_15, gm_n1622, gm_n335);
	nand (gm_n1624, gm_n337, in_27, gm_n158, gm_n1623, gm_n459);
	nor (gm_n1625, gm_n1624, gm_n55);
	and (gm_n1626, gm_n594, gm_n144);
	nand (gm_n1627, gm_n313, in_15, in_11, gm_n1626, gm_n930);
	nor (gm_n1628, gm_n317, gm_n158, in_19, gm_n1627, gm_n360);
	nand (gm_n1629, gm_n182, in_31, gm_n54, gm_n1628, gm_n306);
	nor (gm_n1630, gm_n116, gm_n95, in_8, gm_n599);
	nand (gm_n1631, gm_n302, gm_n58, gm_n62, gm_n1630, gm_n426);
	nor (gm_n1632, gm_n1112, in_27, gm_n158, gm_n1631, gm_n514);
	nand (gm_n1633, gm_n1632, gm_n674, in_31);
	nand (gm_n1634, gm_n396, gm_n264, gm_n124);
	nor (gm_n1635, gm_n236, gm_n73, in_12, gm_n1634, gm_n352);
	nand (gm_n1636, gm_n103, in_24, in_20, gm_n1635, gm_n477);
	nor (gm_n1637, gm_n140, gm_n185, in_28, gm_n1636);
	nor (gm_n1638, gm_n111, gm_n63, gm_n124, gm_n369, gm_n236);
	nand (gm_n1639, gm_n217, in_20, gm_n73, gm_n1638, gm_n521);
	nor (gm_n1640, gm_n226, in_28, gm_n82, gm_n1639, gm_n368);
	nand (gm_n1641, gm_n594, gm_n264, gm_n124);
	or (gm_n1642, gm_n154, in_16, gm_n63, gm_n1641, gm_n188);
	nor (gm_n1643, gm_n187, gm_n82, in_20, gm_n1642, gm_n801);
	nand (gm_n1644, gm_n215, gm_n101, gm_n83, gm_n1643);
	or (gm_n1645, gm_n92, gm_n63, in_8, gm_n1038, gm_n109);
	nor (gm_n1646, gm_n801, gm_n76, gm_n73, gm_n1645, gm_n412);
	nand (gm_n1647, gm_n367, gm_n83, in_24, gm_n1646, gm_n496);
	nor (gm_n1648, gm_n321, in_15, in_11, gm_n991, gm_n619);
	nand (gm_n1649, gm_n334, in_23, in_19, gm_n1648, gm_n359);
	nor (gm_n1650, gm_n57, in_31, gm_n54, gm_n1649, gm_n977);
	nand (gm_n1651, gm_n730, gm_n502, gm_n218);
	nor (gm_n1652, gm_n122, gm_n62, gm_n61, gm_n1651, gm_n991);
	nand (gm_n1653, gm_n60, gm_n158, gm_n58, gm_n1652, gm_n513);
	nor (gm_n1654, gm_n423, in_31, in_27, gm_n1653);
	nor (gm_n1655, gm_n249, in_12, gm_n124, gm_n1034, gm_n111);
	nand (gm_n1656, gm_n107, gm_n76, gm_n73, gm_n1655, gm_n205);
	nor (gm_n1657, gm_n248, gm_n83, gm_n82, gm_n1656, gm_n195);
	nand (gm_n1658, gm_n128, gm_n218, in_11, gm_n698, gm_n300);
	nor (gm_n1659, gm_n796, in_19, in_15, gm_n1658, gm_n317);
	nand (gm_n1660, gm_n60, in_27, in_23, gm_n1659, gm_n337);
	nor (gm_n1661, gm_n1660, gm_n55);
	nor (gm_n1662, gm_n669, gm_n62, in_11, gm_n395, gm_n146);
	nand (gm_n1663, gm_n74, in_23, gm_n58, gm_n1662, gm_n130);
	nor (gm_n1664, gm_n512, in_31, in_27, gm_n1663, gm_n423);
	nor (gm_n1665, gm_n1657, gm_n1654, gm_n1650, gm_n1664, gm_n1661);
	nor (gm_n1666, gm_n374, in_12, in_8, gm_n1038, gm_n237);
	nand (gm_n1667, gm_n107, gm_n76, gm_n73, gm_n1666, gm_n205);
	nor (gm_n1668, gm_n85, in_28, in_24, gm_n1667, gm_n479);
	nor (gm_n1669, gm_n425, gm_n62, in_11, gm_n822, gm_n664);
	nand (gm_n1670, gm_n121, in_23, in_19, gm_n1669, gm_n296);
	nor (gm_n1671, gm_n183, in_31, gm_n54, gm_n1670, gm_n675);
	nor (gm_n1672, gm_n553, gm_n73, in_12, gm_n1296, gm_n237);
	nand (gm_n1673, gm_n164, gm_n82, gm_n76, gm_n1672, gm_n217);
	nor (gm_n1674, gm_n248, gm_n138, gm_n83, gm_n1673);
	nor (gm_n1675, gm_n1674, gm_n1671, gm_n1668);
	and (gm_n1676, in_6, gm_n70, gm_n113, gm_n543, gm_n151);
	nand (gm_n1677, gm_n175, in_12, gm_n61, gm_n1676, gm_n300);
	nor (gm_n1678, gm_n157, in_21, gm_n105, gm_n1677, gm_n767);
	nor (gm_n1679, in_28, gm_n54, gm_n59);
	nand (gm_n1680, gm_n539, gm_n80, gm_n133, gm_n1679, gm_n1678);
	nor (gm_n1681, gm_n1680, gm_n55, in_30);
	nand (gm_n1682, gm_n127, in_12, gm_n124, gm_n502, gm_n256);
	nor (gm_n1683, gm_n236, in_20, in_16, gm_n1682, gm_n476);
	nand (gm_n1684, gm_n102, gm_n83, gm_n82, gm_n1683, gm_n227);
	nor (gm_n1685, gm_n1684, gm_n684);
	nand (gm_n1686, gm_n402, gm_n144, in_8);
	nor (gm_n1687, gm_n249, in_16, in_12, gm_n1686, gm_n282);
	nand (gm_n1688, gm_n107, gm_n82, in_20, gm_n1687, gm_n255);
	nor (gm_n1689, gm_n262, gm_n185, gm_n83, gm_n1688);
	nor (gm_n1690, gm_n1689, gm_n1685, gm_n1681);
	nand (gm_n1691, gm_n1665, gm_n1647, gm_n1644, gm_n1690, gm_n1675);
	and (gm_n1692, gm_n649, in_17, in_13, gm_n1125, gm_n733);
	and (gm_n1693, gm_n540, in_25, in_21, gm_n1692, gm_n1180);
	nand (gm_n1694, gm_n55, gm_n100, gm_n80, gm_n1693);
	nand (gm_n1695, gm_n797, in_15, in_11, gm_n622, gm_n544);
	nor (gm_n1696, gm_n1225, in_23, in_19, gm_n1695, gm_n613);
	nand (gm_n1697, gm_n182, gm_n55, gm_n54, gm_n1696, gm_n674);
	nor (gm_n1698, gm_n93, in_12, gm_n124, gm_n168, gm_n154);
	nand (gm_n1699, gm_n141, gm_n76, in_16, gm_n1698, gm_n207);
	nor (gm_n1700, gm_n104, in_28, gm_n82, gm_n1699, gm_n140);
	nand (gm_n1701, gm_n1700, gm_n196);
	nand (gm_n1702, gm_n1701, gm_n1697, gm_n1694);
	or (gm_n1703, gm_n92, in_16, gm_n63, gm_n1168, gm_n553);
	nor (gm_n1704, gm_n520, in_24, in_20, gm_n1703, gm_n412);
	nand (gm_n1705, gm_n196, gm_n139, in_28, gm_n1704);
	nor (gm_n1706, gm_n277, gm_n152, in_8);
	nand (gm_n1707, gm_n199, gm_n74, in_15, gm_n1706, gm_n622);
	nor (gm_n1708, gm_n183, in_23, in_19, gm_n1707, gm_n514);
	nand (gm_n1709, gm_n306, in_31, gm_n54, gm_n1708);
	and (gm_n1710, gm_n115, gm_n70, gm_n113, gm_n543, in_7);
	nand (gm_n1711, gm_n126, gm_n62, in_11, gm_n1710, gm_n622);
	nor (gm_n1712, gm_n303, in_23, gm_n58, gm_n1711, gm_n317);
	nand (gm_n1713, gm_n134, in_31, gm_n54, gm_n1712, gm_n674);
	nand (gm_n1714, gm_n1713, gm_n1709, gm_n1705);
	nor (gm_n1715, gm_n1691, gm_n1640, gm_n1637, gm_n1714, gm_n1702);
	nor (gm_n1716, gm_n374, gm_n63, gm_n124, gm_n600, gm_n282);
	nand (gm_n1717, gm_n192, gm_n76, gm_n73, gm_n1716, gm_n477);
	nor (gm_n1718, gm_n85, in_28, gm_n82, gm_n1717, gm_n479);
	nand (gm_n1719, gm_n588, gm_n218, gm_n124);
	nor (gm_n1720, gm_n92, in_16, gm_n63, gm_n1719, gm_n177);
	nand (gm_n1721, gm_n164, in_24, in_20, gm_n1720, gm_n205);
	nor (gm_n1722, gm_n262, gm_n226, gm_n83, gm_n1721);
	nand (gm_n1723, gm_n703, gm_n71);
	nor (gm_n1724, gm_n363, gm_n62, gm_n61, gm_n1723, gm_n664);
	nand (gm_n1725, gm_n392, in_23, in_19, gm_n1724, gm_n513);
	nor (gm_n1726, gm_n183, gm_n55, gm_n54, gm_n1725, gm_n838);
	nor (gm_n1727, gm_n1726, gm_n1722, gm_n1718);
	nor (gm_n1728, gm_n92, gm_n63, in_8, gm_n739, gm_n143);
	nand (gm_n1729, gm_n217, gm_n76, in_16, gm_n1728, gm_n235);
	nor (gm_n1730, gm_n224, gm_n83, gm_n82, gm_n1729, gm_n684);
	and (gm_n1731, in_8, in_4, gm_n68, gm_n145, gm_n144);
	and (gm_n1732, gm_n110, gm_n73, in_12, gm_n1731, gm_n142);
	nand (gm_n1733, gm_n164, in_24, in_20, gm_n1732, gm_n217);
	nor (gm_n1734, gm_n214, gm_n140, in_28, gm_n1733);
	nor (gm_n1735, gm_n92, in_16, in_12, gm_n1019, gm_n236);
	nand (gm_n1736, gm_n90, in_24, in_20, gm_n1735, gm_n263);
	nor (gm_n1737, gm_n138, gm_n224, in_28, gm_n1736);
	nor (gm_n1738, gm_n1737, gm_n1734, gm_n1730);
	nand (gm_n1739, gm_n1715, gm_n1633, gm_n1629, gm_n1738, gm_n1727);
	and (gm_n1740, gm_n731, gm_n127, in_8);
	nand (gm_n1741, gm_n199, in_16, gm_n63, gm_n1740, gm_n207);
	nor (gm_n1742, gm_n165, in_24, in_20, gm_n1741, gm_n801);
	nand (gm_n1743, gm_n213, gm_n84, gm_n83, gm_n1742);
	and (gm_n1744, gm_n219, gm_n153, in_8, gm_n264);
	nand (gm_n1745, gm_n302, in_19, gm_n62, gm_n1744, gm_n1226);
	nor (gm_n1746, gm_n297, gm_n54, gm_n158, gm_n1745, gm_n1200);
	nand (gm_n1747, gm_n1746, gm_n306, in_31);
	and (gm_n1748, gm_n243, gm_n218, gm_n61, gm_n426, gm_n300);
	nand (gm_n1749, gm_n121, in_19, in_15, gm_n1748, gm_n513);
	nor (gm_n1750, gm_n612, in_27, gm_n158, gm_n1749, gm_n458);
	nand (gm_n1751, gm_n1750, in_31);
	nand (gm_n1752, gm_n1751, gm_n1747, gm_n1743);
	nand (gm_n1753, gm_n110, gm_n73, in_12, gm_n1331, gm_n207);
	nor (gm_n1754, gm_n165, in_24, gm_n76, gm_n1753, gm_n566);
	nand (gm_n1755, gm_n215, gm_n137, in_28, gm_n1754);
	and (gm_n1756, gm_n110, gm_n63, in_8, gm_n703, gm_n189);
	nand (gm_n1757, gm_n207, gm_n76, in_16, gm_n1756, gm_n270);
	nor (gm_n1758, gm_n224, in_28, gm_n82, gm_n1757, gm_n206);
	nand (gm_n1759, gm_n1758, gm_n196);
	and (gm_n1760, gm_n515, gm_n289);
	nand (gm_n1761, gm_n394, gm_n62, in_11, gm_n1760, gm_n931);
	nor (gm_n1762, gm_n796, in_23, gm_n58, gm_n1761, gm_n452);
	nand (gm_n1763, gm_n134, gm_n55, in_27, gm_n1762, gm_n511);
	nand (gm_n1764, gm_n1763, gm_n1759, gm_n1755);
	nor (gm_n1765, gm_n1739, gm_n1625, gm_n1621, gm_n1764, gm_n1752);
	and (gm_n1766, gm_n150, in_16, in_12, gm_n1355, gm_n153);
	nand (gm_n1767, gm_n263, in_24, gm_n76, gm_n1766, gm_n270);
	nor (gm_n1768, gm_n226, gm_n85, in_28, gm_n1767);
	nor (gm_n1769, gm_n109, gm_n73, in_12, gm_n1296, gm_n237);
	nand (gm_n1770, gm_n141, in_24, gm_n76, gm_n1769, gm_n217);
	nor (gm_n1771, gm_n226, gm_n216, in_28, gm_n1770);
	nand (gm_n1772, gm_n402, gm_n515, in_8);
	nor (gm_n1773, gm_n143, gm_n73, gm_n63, gm_n1772, gm_n599);
	nand (gm_n1774, gm_n227, in_24, in_20, gm_n1773, gm_n521);
	nor (gm_n1775, gm_n368, gm_n226, gm_n83, gm_n1774);
	nor (gm_n1776, gm_n1775, gm_n1771, gm_n1768);
	nand (gm_n1777, gm_n90, in_24, gm_n76, gm_n922, gm_n263);
	nor (gm_n1778, gm_n368, gm_n214, in_28, gm_n1777);
	nand (gm_n1779, gm_n264, gm_n63, gm_n124, gm_n311, gm_n340);
	nor (gm_n1780, gm_n249, gm_n76, in_16, gm_n1779, gm_n476);
	nand (gm_n1781, gm_n139, gm_n83, in_24, gm_n1780, gm_n205);
	nor (gm_n1782, gm_n1781, gm_n234);
	nor (gm_n1783, gm_n670, gm_n62, gm_n61, gm_n1209, gm_n425);
	nand (gm_n1784, gm_n173, in_23, in_19, gm_n1783, gm_n174);
	nor (gm_n1785, gm_n423, in_31, gm_n54, gm_n1784, gm_n458);
	nor (gm_n1786, gm_n1785, gm_n1782, gm_n1778);
	nand (gm_n1787, gm_n1765, gm_n1617, gm_n1612, gm_n1786, gm_n1776);
	nand (gm_n1788, gm_n200, gm_n73, in_12, gm_n516, gm_n242);
	nor (gm_n1789, gm_n187, gm_n82, gm_n76, gm_n1788, gm_n520);
	nand (gm_n1790, gm_n496, gm_n186, gm_n83, gm_n1789);
	nor (gm_n1791, gm_n383, gm_n114);
	nand (gm_n1792, gm_n730, in_15, gm_n61, gm_n1791, gm_n1226);
	nor (gm_n1793, gm_n452, in_23, gm_n58, gm_n1792, gm_n456);
	nand (gm_n1794, gm_n134, in_31, in_27, gm_n1793, gm_n438);
	nand (gm_n1795, gm_n283, gm_n71, gm_n124);
	or (gm_n1796, gm_n236, gm_n73, gm_n63, gm_n1795, gm_n599);
	nor (gm_n1797, gm_n89, gm_n82, in_20, gm_n1796, gm_n197);
	nand (gm_n1798, gm_n496, gm_n139, in_28, gm_n1797);
	nand (gm_n1799, gm_n1798, gm_n1794, gm_n1790);
	nand (gm_n1800, gm_n144, in_12, gm_n124, gm_n242, gm_n208);
	nor (gm_n1801, gm_n187, gm_n76, in_16, gm_n1800, gm_n188);
	nand (gm_n1802, gm_n103, gm_n83, in_24, gm_n1801, gm_n186);
	nor (gm_n1803, gm_n1802, gm_n479);
	nor (out_6, gm_n1799, gm_n1787, gm_n1609, gm_n1803);
	nand (gm_n1805, gm_n594, gm_n218);
	nor (gm_n1806, gm_n143, gm_n63, in_8, gm_n1805, gm_n288);
	nand (gm_n1807, gm_n88, in_20, in_16, gm_n1806, gm_n270);
	nor (gm_n1808, gm_n140, gm_n83, gm_n82, gm_n1807, gm_n195);
	nand (gm_n1809, gm_n91, in_16, in_12, gm_n230, gm_n199);
	nor (gm_n1810, gm_n197, gm_n82, in_20, gm_n1809, gm_n104);
	nand (gm_n1811, gm_n213, gm_n139, in_28, gm_n1810);
	nand (gm_n1812, gm_n446, in_16, in_12, gm_n1363, gm_n228);
	nor (gm_n1813, gm_n197, gm_n82, gm_n76, gm_n1812, gm_n801);
	nand (gm_n1814, gm_n196, gm_n186, in_28, gm_n1813);
	nor (gm_n1815, gm_n432, gm_n62, gm_n61, gm_n1272, gm_n395);
	nand (gm_n1816, gm_n513, in_23, gm_n58, gm_n1815, gm_n1042);
	nor (gm_n1817, gm_n1200, gm_n55, gm_n54, gm_n1816, gm_n618);
	nand (gm_n1818, gm_n289, gm_n264, in_11, gm_n394, gm_n313);
	nor (gm_n1819, gm_n431, gm_n58, in_15, gm_n1818, gm_n613);
	nand (gm_n1820, gm_n309, gm_n54, in_23, gm_n1819, gm_n438);
	nor (gm_n1821, gm_n1820, gm_n55);
	nand (gm_n1822, gm_n65, gm_n58, gm_n62, gm_n1744, gm_n174);
	nor (gm_n1823, gm_n452, in_27, in_23, gm_n1822, gm_n183);
	nand (gm_n1824, gm_n1823, gm_n56, gm_n55);
	nor (gm_n1825, gm_n178, in_12, in_8, gm_n345, gm_n237);
	nand (gm_n1826, gm_n90, gm_n76, in_16, gm_n1825, gm_n200);
	nor (gm_n1827, gm_n206, gm_n83, in_24, gm_n1826, gm_n368);
	nand (gm_n1828, gm_n1827, gm_n81);
	nand (gm_n1829, gm_n153, in_12, gm_n124, gm_n703, gm_n310);
	nor (gm_n1830, gm_n177, gm_n76, gm_n73, gm_n1829, gm_n476);
	nand (gm_n1831, gm_n186, in_28, in_24, gm_n1830, gm_n192);
	nor (gm_n1832, gm_n1831, gm_n226);
	nor (gm_n1833, gm_n553, gm_n63, in_8, gm_n503, gm_n288);
	nand (gm_n1834, gm_n88, gm_n76, in_16, gm_n1833, gm_n90);
	nor (gm_n1835, gm_n224, gm_n83, in_24, gm_n1834, gm_n479);
	nor (gm_n1836, gm_n151, gm_n115, gm_n70, gm_n229, in_8);
	nand (gm_n1837, gm_n176, in_16, gm_n63, gm_n1836, gm_n256);
	nor (gm_n1838, gm_n197, in_24, in_20, gm_n1837, gm_n630);
	nand (gm_n1839, gm_n225, gm_n84, gm_n83, gm_n1838);
	nor (gm_n1840, in_16, gm_n62, gm_n64);
	nor (gm_n1841, gm_n345, gm_n198, gm_n124, gm_n548);
	nor (gm_n1842, gm_n63, gm_n61, in_10);
	and (gm_n1843, gm_n1840, in_17, in_13, gm_n1842, gm_n1841);
	and (gm_n1844, gm_n407, in_25, gm_n86, gm_n1843, gm_n531);
	nand (gm_n1845, gm_n55, gm_n100, in_29, gm_n1844, gm_n735);
	nor (gm_n1846, gm_n109, gm_n63, in_8, gm_n822, gm_n352);
	nand (gm_n1847, gm_n217, in_20, gm_n73, gm_n1846, gm_n235);
	nor (gm_n1848, gm_n138, in_28, in_24, gm_n1847, gm_n140);
	nor (gm_n1849, gm_n599, in_12, gm_n124, gm_n384, gm_n177);
	nand (gm_n1850, gm_n164, in_20, in_16, gm_n1849, gm_n255);
	nor (gm_n1851, gm_n138, gm_n83, in_24, gm_n1850, gm_n774);
	nor (gm_n1852, gm_n154, gm_n63, gm_n124, gm_n1527, gm_n188);
	nand (gm_n1853, gm_n164, gm_n76, in_16, gm_n1852, gm_n192);
	nor (gm_n1854, gm_n138, gm_n83, in_24, gm_n1853, gm_n140);
	nand (gm_n1855, gm_n144, gm_n69);
	nor (gm_n1856, gm_n249, in_12, gm_n124, gm_n1855, gm_n599);
	nand (gm_n1857, gm_n255, in_20, in_16, gm_n1856, gm_n521);
	nor (gm_n1858, gm_n85, gm_n83, gm_n82, gm_n1857, gm_n479);
	nand (gm_n1859, gm_n71, in_12, gm_n124, gm_n1033, gm_n110);
	nor (gm_n1860, gm_n249, in_20, gm_n73, gm_n1859, gm_n187);
	nand (gm_n1861, gm_n205, in_28, gm_n82, gm_n1860, gm_n339);
	nor (gm_n1862, gm_n1861, gm_n226);
	nor (gm_n1863, gm_n1854, gm_n1851, gm_n1848, gm_n1862, gm_n1858);
	nor (gm_n1864, gm_n146, gm_n62, in_11, gm_n398, gm_n322);
	nand (gm_n1865, gm_n316, in_23, in_19, gm_n1864, gm_n392);
	nor (gm_n1866, gm_n1112, gm_n55, in_27, gm_n1865, gm_n423);
	nor (gm_n1867, gm_n670, in_15, in_11, gm_n397, gm_n363);
	nand (gm_n1868, gm_n121, gm_n158, gm_n58, gm_n1867, gm_n173);
	nor (gm_n1869, gm_n458, in_31, gm_n54, gm_n1868, gm_n675);
	nand (gm_n1870, gm_n144, gm_n63, gm_n124, gm_n775, gm_n242);
	nor (gm_n1871, gm_n109, in_20, in_16, gm_n1870, gm_n522);
	nand (gm_n1872, gm_n186, in_28, gm_n82, gm_n1871, gm_n263);
	nor (gm_n1873, gm_n1872, gm_n226);
	nor (gm_n1874, gm_n1873, gm_n1869, gm_n1866);
	nor (gm_n1875, gm_n669, gm_n62, gm_n61, gm_n600, gm_n670);
	nand (gm_n1876, gm_n74, gm_n158, in_19, gm_n1875, gm_n334);
	nor (gm_n1877, gm_n422, gm_n55, in_27, gm_n1876, gm_n423);
	nor (gm_n1878, gm_n109, gm_n73, gm_n63, gm_n290, gm_n154);
	nand (gm_n1879, gm_n164, in_24, gm_n76, gm_n1878, gm_n227);
	nor (gm_n1880, gm_n262, gm_n234, in_28, gm_n1879);
	or (gm_n1881, gm_n383, gm_n229, in_8);
	nor (gm_n1882, gm_n177, in_16, in_12, gm_n1881, gm_n282);
	nand (gm_n1883, gm_n235, in_24, in_20, gm_n1882, gm_n255);
	nor (gm_n1884, gm_n262, gm_n226, in_28, gm_n1883);
	nor (gm_n1885, gm_n1884, gm_n1880, gm_n1877);
	nand (gm_n1886, gm_n1863, gm_n1845, gm_n1839, gm_n1885, gm_n1874);
	and (gm_n1887, gm_n515, gm_n243, gm_n124);
	nand (gm_n1888, gm_n153, in_16, in_12, gm_n1887, gm_n176);
	nor (gm_n1889, gm_n197, in_24, in_20, gm_n1888, gm_n520);
	nand (gm_n1890, gm_n225, gm_n139, in_28, gm_n1889);
	nor (gm_n1891, in_21, in_20);
	nand (gm_n1892, gm_n256, in_12, gm_n124, gm_n310, gm_n283);
	nor (gm_n1893, gm_n1892, gm_n64, gm_n175);
	nand (gm_n1894, gm_n486, in_19, gm_n106, gm_n1893, gm_n1891);
	nand (gm_n1895, gm_n133, gm_n82, in_23);
	nor (gm_n1896, gm_n1894, in_26, in_22, gm_n1895);
	nor (gm_n1897, in_29, gm_n83, in_27);
	nand (gm_n1898, gm_n1896, gm_n55, gm_n100, gm_n1897);
	and (gm_n1899, gm_n151, in_6, gm_n70, gm_n361);
	nand (gm_n1900, gm_n142, in_12, gm_n124, gm_n1899, gm_n242);
	nor (gm_n1901, gm_n89, gm_n76, in_16, gm_n1900, gm_n108);
	nand (gm_n1902, gm_n186, in_28, gm_n82, gm_n1901, gm_n196);
	nand (gm_n1903, gm_n1902, gm_n1898, gm_n1890);
	nor (gm_n1904, gm_n535, in_8, in_7);
	nand (gm_n1905, gm_n359, gm_n242, gm_n62, gm_n1904, gm_n931);
	nor (gm_n1906, gm_n1225, in_23, gm_n58, gm_n1905, gm_n422);
	nand (gm_n1907, gm_n308, in_31, gm_n54, gm_n1906);
	nand (gm_n1908, gm_n110, in_16, gm_n63, gm_n562, gm_n176);
	nor (gm_n1909, gm_n108, in_24, gm_n76, gm_n1908, gm_n411);
	nand (gm_n1910, gm_n102, gm_n81, in_28, gm_n1909);
	or (gm_n1911, gm_n599, gm_n73, in_12, gm_n1541, gm_n188);
	nor (gm_n1912, gm_n89, in_24, gm_n76, gm_n1911, gm_n412);
	nand (gm_n1913, gm_n215, gm_n196, in_28, gm_n1912);
	nand (gm_n1914, gm_n1913, gm_n1910, gm_n1907);
	nor (gm_n1915, gm_n1886, gm_n1835, gm_n1832, gm_n1914, gm_n1903);
	nor (gm_n1916, gm_n109, in_16, gm_n63, gm_n353, gm_n154);
	nand (gm_n1917, gm_n107, in_24, gm_n76, gm_n1916, gm_n227);
	nor (gm_n1918, gm_n774, gm_n214, in_28, gm_n1917);
	nand (gm_n1919, gm_n167, in_12, gm_n124, gm_n588, gm_n515);
	nor (gm_n1920, gm_n108, in_20, in_16, gm_n1919, gm_n188);
	nand (gm_n1921, gm_n227, gm_n83, gm_n82, gm_n1920, gm_n466);
	nor (gm_n1922, gm_n1921, gm_n214);
	nor (gm_n1923, gm_n177, in_16, gm_n63, gm_n1795, gm_n282);
	nand (gm_n1924, gm_n164, gm_n82, gm_n76, gm_n1923, gm_n192);
	nor (gm_n1925, gm_n479, gm_n368, gm_n83, gm_n1924);
	nor (gm_n1926, gm_n1925, gm_n1922, gm_n1918);
	nor (gm_n1927, gm_n374, in_16, gm_n63, gm_n1117, gm_n282);
	nand (gm_n1928, gm_n107, gm_n82, gm_n76, gm_n1927, gm_n192);
	nor (gm_n1929, gm_n226, gm_n248, in_28, gm_n1928);
	and (gm_n1930, gm_n153, gm_n73, in_12, gm_n981, gm_n446);
	nand (gm_n1931, gm_n103, in_24, in_20, gm_n1930, gm_n164);
	nor (gm_n1932, gm_n262, gm_n226, gm_n83, gm_n1931);
	and (gm_n1933, gm_n797, in_15, gm_n61, gm_n544, gm_n931);
	nand (gm_n1934, gm_n130, gm_n158, in_19, gm_n1933, gm_n302);
	nor (gm_n1935, gm_n512, in_31, in_27, gm_n1934, gm_n612);
	nor (gm_n1936, gm_n1935, gm_n1932, gm_n1929);
	nand (gm_n1937, gm_n1915, gm_n1828, gm_n1824, gm_n1936, gm_n1926);
	and (gm_n1938, gm_n620, gm_n515);
	nand (gm_n1939, gm_n126, gm_n62, in_11, gm_n1938, gm_n1226);
	nor (gm_n1940, gm_n297, in_23, in_19, gm_n1939, gm_n393);
	nand (gm_n1941, gm_n60, gm_n55, in_27, gm_n1940, gm_n674);
	and (gm_n1942, gm_n283, gm_n71, in_11, gm_n931, gm_n394);
	nand (gm_n1943, gm_n296, gm_n58, gm_n62, gm_n1942, gm_n302);
	nor (gm_n1944, gm_n458, in_27, in_23, gm_n1943, gm_n675);
	nand (gm_n1945, gm_n1944, gm_n55);
	and (gm_n1946, gm_n396, gm_n144);
	nand (gm_n1947, gm_n200, in_12, gm_n124, gm_n1946, gm_n228);
	nor (gm_n1948, gm_n411, gm_n76, gm_n73, gm_n1947, gm_n412);
	nand (gm_n1949, gm_n339, in_28, gm_n82, gm_n1948, gm_n629);
	nand (gm_n1950, gm_n1949, gm_n1945, gm_n1941);
	or (gm_n1951, gm_n177, in_16, in_12, gm_n375, gm_n288);
	nor (gm_n1952, gm_n165, gm_n82, in_20, gm_n1951, gm_n566);
	nand (gm_n1953, gm_n496, gm_n466, gm_n83, gm_n1952);
	nand (gm_n1954, gm_n65, gm_n62, gm_n61, gm_n1195, gm_n730);
	nor (gm_n1955, gm_n122, in_23, gm_n58, gm_n1954, gm_n317);
	nand (gm_n1956, gm_n182, gm_n55, gm_n54, gm_n1955, gm_n674);
	nand (gm_n1957, gm_n150, in_16, in_12, gm_n754, gm_n228);
	nor (gm_n1958, gm_n463, in_24, gm_n76, gm_n1957, gm_n630);
	nand (gm_n1959, gm_n213, gm_n186, in_28, gm_n1958);
	nand (gm_n1960, gm_n1959, gm_n1956, gm_n1953);
	nor (gm_n1961, gm_n1937, gm_n1821, gm_n1817, gm_n1960, gm_n1950);
	nor (gm_n1962, gm_n670, in_15, in_11, gm_n584, gm_n425);
	nand (gm_n1963, gm_n296, gm_n158, in_19, gm_n1962, gm_n302);
	nor (gm_n1964, gm_n512, in_31, gm_n54, gm_n1963, gm_n618);
	nand (gm_n1965, gm_n242, gm_n189, gm_n124, gm_n502);
	nor (gm_n1966, gm_n249, in_16, gm_n63, gm_n1965, gm_n476);
	nand (gm_n1967, gm_n84, gm_n82, gm_n76, gm_n1966, gm_n227);
	nor (gm_n1968, gm_n1967, gm_n479, gm_n83);
	nor (gm_n1969, gm_n433, in_15, gm_n61, gm_n1252, gm_n363);
	nand (gm_n1970, gm_n173, in_23, gm_n58, gm_n1969, gm_n455);
	nor (gm_n1971, gm_n57, gm_n55, gm_n54, gm_n1970, gm_n183);
	nor (gm_n1972, gm_n1971, gm_n1968, gm_n1964);
	nor (gm_n1973, gm_n249, gm_n73, gm_n63, gm_n1287, gm_n282);
	nand (gm_n1974, gm_n263, in_24, in_20, gm_n1973, gm_n270);
	nor (gm_n1975, gm_n479, gm_n224, gm_n83, gm_n1974);
	nor (gm_n1976, gm_n393, gm_n58, gm_n62, gm_n925, gm_n398);
	nand (gm_n1977, gm_n130, gm_n54, gm_n158, gm_n1976, gm_n391);
	nor (gm_n1978, gm_n1977, gm_n357, gm_n55);
	nand (gm_n1979, gm_n151, in_6, in_5, gm_n361, gm_n124);
	nor (gm_n1980, gm_n188, gm_n73, gm_n63, gm_n1979, gm_n237);
	nand (gm_n1981, gm_n107, gm_n82, gm_n76, gm_n1980, gm_n217);
	nor (gm_n1982, gm_n226, gm_n216, gm_n83, gm_n1981);
	nor (gm_n1983, gm_n1982, gm_n1978, gm_n1975);
	nand (gm_n1984, gm_n1961, gm_n1814, gm_n1811, gm_n1983, gm_n1972);
	nand (gm_n1985, gm_n91, in_16, in_12, gm_n784, gm_n228);
	nor (gm_n1986, gm_n187, in_24, gm_n76, gm_n1985, gm_n801);
	nand (gm_n1987, gm_n102, gm_n101, in_28, gm_n1986);
	nor (gm_n1988, in_9, in_8, in_7);
	nand (gm_n1989, in_10, in_6, in_5, gm_n1988, gm_n283);
	nor (gm_n1990, gm_n1989, gm_n61);
	nand (gm_n1991, gm_n121, in_19, in_15, gm_n1990, gm_n123);
	nor (gm_n1992, gm_n422, gm_n54, gm_n158, gm_n1991, gm_n514);
	nand (gm_n1993, gm_n1992, gm_n511, gm_n55);
	and (gm_n1994, gm_n588, gm_n264, in_8);
	nand (gm_n1995, gm_n200, in_16, gm_n63, gm_n1994, gm_n340);
	nor (gm_n1996, gm_n206, gm_n82, in_20, gm_n1995, gm_n522);
	nand (gm_n1997, gm_n215, gm_n213, gm_n83, gm_n1996);
	nand (gm_n1998, gm_n1997, gm_n1993, gm_n1987);
	and (gm_n1999, gm_n515, gm_n242, gm_n124, gm_n703);
	and (gm_n2000, gm_n65, gm_n58, gm_n62, gm_n1999, gm_n392);
	nand (gm_n2001, gm_n130, in_27, in_23, gm_n2000, gm_n182);
	nor (gm_n2002, gm_n2001, gm_n357, gm_n55);
	nor (out_7, gm_n1998, gm_n1984, gm_n1808, gm_n2002);
	nor (gm_n2004, gm_n249, gm_n73, in_12, gm_n896, gm_n111);
	nand (gm_n2005, gm_n217, in_24, in_20, gm_n2004, gm_n235);
	nor (gm_n2006, gm_n262, gm_n226, gm_n83, gm_n2005);
	nor (gm_n2007, in_12, in_11, gm_n66);
	nand (gm_n2008, gm_n533, gm_n105, gm_n175, gm_n2007, gm_n1841);
	nand (gm_n2009, in_24, gm_n158, gm_n87);
	nor (gm_n2010, gm_n157, in_25, in_21, gm_n2009, gm_n2008);
	nand (gm_n2011, gm_n55, in_30, gm_n80, gm_n2010, gm_n1679);
	and (gm_n2012, gm_n588, gm_n127, gm_n124);
	nand (gm_n2013, gm_n200, in_16, in_12, gm_n2012, gm_n153);
	nor (gm_n2014, gm_n801, gm_n82, gm_n76, gm_n2013, gm_n412);
	nand (gm_n2015, gm_n339, gm_n137, gm_n83, gm_n2014);
	nor (gm_n2016, gm_n177, gm_n73, in_12, gm_n1965, gm_n476);
	nand (gm_n2017, gm_n263, in_24, in_20, gm_n2016, gm_n367);
	nor (gm_n2018, gm_n2017, gm_n185, gm_n83);
	and (gm_n2019, gm_n930, in_15, in_11, gm_n1133, gm_n426);
	nand (gm_n2020, gm_n174, gm_n158, gm_n58, gm_n2019, gm_n358);
	nor (gm_n2021, gm_n512, in_31, gm_n54, gm_n2020, gm_n618);
	and (gm_n2022, gm_n127, gm_n69);
	nand (gm_n2023, gm_n797, in_15, in_11, gm_n426, gm_n2022);
	nor (gm_n2024, gm_n796, gm_n158, gm_n58, gm_n2023, gm_n131);
	nand (gm_n2025, gm_n459, gm_n55, gm_n54, gm_n2024, gm_n511);
	or (gm_n2026, gm_n236, in_16, in_12, gm_n631, gm_n352);
	nor (gm_n2027, gm_n463, gm_n82, gm_n76, gm_n2026, gm_n630);
	nand (gm_n2028, gm_n225, gm_n84, gm_n83, gm_n2027);
	nor (gm_n2029, gm_n553, in_16, gm_n63, gm_n1541, gm_n154);
	nand (gm_n2030, gm_n164, gm_n82, gm_n76, gm_n2029, gm_n227);
	nor (gm_n2031, gm_n479, gm_n224, in_28, gm_n2030);
	nand (gm_n2032, gm_n775, gm_n71, in_8);
	nor (gm_n2033, gm_n111, in_16, in_12, gm_n2032, gm_n143);
	nand (gm_n2034, gm_n90, in_24, gm_n76, gm_n2033, gm_n255);
	nor (gm_n2035, gm_n262, gm_n195, in_28, gm_n2034);
	nand (gm_n2036, gm_n446, gm_n73, gm_n63, gm_n1150, gm_n228);
	nor (gm_n2037, gm_n566, in_24, in_20, gm_n2036, gm_n522);
	nand (gm_n2038, gm_n225, gm_n84, gm_n83, gm_n2037);
	nor (gm_n2039, gm_n469, gm_n383, gm_n124);
	nand (gm_n2040, gm_n199, in_16, in_12, gm_n2039, gm_n176);
	nor (gm_n2041, gm_n411, gm_n82, gm_n76, gm_n2040, gm_n412);
	nand (gm_n2042, gm_n367, gm_n137, gm_n83, gm_n2041);
	nor (gm_n2043, gm_n109, gm_n73, in_12, gm_n1046, gm_n282);
	nand (gm_n2044, gm_n88, in_24, in_20, gm_n2043, gm_n477);
	nor (gm_n2045, gm_n195, gm_n224, gm_n83, gm_n2044);
	nand (gm_n2046, gm_n453, gm_n515, in_8);
	nor (gm_n2047, gm_n553, gm_n73, gm_n63, gm_n2046, gm_n237);
	nand (gm_n2048, gm_n88, gm_n82, gm_n76, gm_n2047, gm_n90);
	nor (gm_n2049, gm_n214, gm_n224, in_28, gm_n2048);
	nor (gm_n2050, gm_n393, gm_n58, gm_n62, gm_n925, gm_n623);
	nand (gm_n2051, gm_n173, gm_n54, gm_n158, gm_n2050, gm_n657);
	nor (gm_n2052, gm_n2051, gm_n618, gm_n55);
	and (gm_n2053, gm_n110, gm_n63, in_8, gm_n1400, gm_n166);
	nand (gm_n2054, gm_n107, in_20, in_16, gm_n2053, gm_n255);
	nor (gm_n2055, gm_n248, gm_n83, in_24, gm_n2054, gm_n195);
	nand (gm_n2056, gm_n228, gm_n218, gm_n124, gm_n402);
	nor (gm_n2057, gm_n360, in_19, gm_n62, gm_n2056, gm_n623);
	nand (gm_n2058, gm_n130, in_27, gm_n158, gm_n2057, gm_n459);
	nor (gm_n2059, gm_n2058, gm_n423, gm_n55);
	nor (gm_n2060, gm_n2052, gm_n2049, gm_n2045, gm_n2059, gm_n2055);
	nor (gm_n2061, gm_n143, gm_n63, in_11, gm_n758, gm_n670);
	nand (gm_n2062, gm_n141, in_20, gm_n73, gm_n2061, gm_n217);
	nor (gm_n2063, gm_n224, in_28, in_24, gm_n2062, gm_n684);
	nor (gm_n2064, gm_n154, in_16, gm_n63, gm_n1359, gm_n236);
	nand (gm_n2065, gm_n88, gm_n82, gm_n76, gm_n2064, gm_n477);
	nor (gm_n2066, gm_n684, gm_n248, gm_n83, gm_n2065);
	nand (gm_n2067, gm_n296, in_23, in_19, gm_n1139, gm_n1042);
	nor (gm_n2068, gm_n423, gm_n55, in_27, gm_n2067, gm_n458);
	nor (gm_n2069, gm_n2068, gm_n2066, gm_n2063);
	nand (gm_n2070, gm_n310, gm_n69, in_8);
	nor (gm_n2071, gm_n154, gm_n669, in_15, gm_n2070, gm_n613);
	nand (gm_n2072, gm_n305, gm_n158, in_19, gm_n2071, gm_n513);
	nor (gm_n2073, gm_n423, gm_n55, gm_n54, gm_n2072);
	nand (gm_n2074, gm_n402, gm_n71);
	nor (gm_n2075, gm_n395, in_15, in_11, gm_n2074, gm_n398);
	nand (gm_n2076, gm_n77, in_23, gm_n58, gm_n2075, gm_n359);
	nor (gm_n2077, gm_n838, in_31, gm_n54, gm_n2076, gm_n977);
	nor (gm_n2078, gm_n664, gm_n62, in_11, gm_n1805, gm_n991);
	nand (gm_n2079, gm_n296, gm_n158, in_19, gm_n2078, gm_n302);
	nor (gm_n2080, gm_n1200, gm_n55, in_27, gm_n2079, gm_n437);
	nor (gm_n2081, gm_n2080, gm_n2077, gm_n2073);
	nand (gm_n2082, gm_n2060, gm_n2042, gm_n2038, gm_n2081, gm_n2069);
	nand (gm_n2083, gm_n91, gm_n76, gm_n73, gm_n477, gm_n244);
	nor (gm_n2084, gm_n206, in_28, gm_n82, gm_n2083, gm_n774);
	nand (gm_n2085, gm_n2084, gm_n496);
	nand (gm_n2086, gm_n150, in_16, in_12, gm_n1887, gm_n242);
	nor (gm_n2087, gm_n165, gm_n82, gm_n76, gm_n2086, gm_n630);
	nand (gm_n2088, gm_n102, gm_n101, gm_n83, gm_n2087);
	nand (gm_n2089, gm_n931, gm_n62, in_11, gm_n1676, gm_n424);
	nor (gm_n2090, gm_n796, gm_n158, gm_n58, gm_n2089, gm_n317);
	nand (gm_n2091, gm_n337, gm_n55, gm_n54, gm_n2090, gm_n459);
	nand (gm_n2092, gm_n2091, gm_n2088, gm_n2085);
	nand (gm_n2093, gm_n797, in_15, gm_n61, gm_n1312, gm_n426);
	nor (gm_n2094, gm_n796, gm_n158, in_19, gm_n2093, gm_n317);
	nand (gm_n2095, gm_n391, in_31, in_27, gm_n2094, gm_n674);
	and (gm_n2096, gm_n588, gm_n71, in_8);
	nand (gm_n2097, gm_n150, in_16, in_12, gm_n2096, gm_n256);
	nor (gm_n2098, gm_n104, in_24, gm_n76, gm_n2097, gm_n165);
	nand (gm_n2099, gm_n186, gm_n137, gm_n83, gm_n2098);
	or (gm_n2100, gm_n432, in_15, gm_n61, gm_n758, gm_n125);
	nor (gm_n2101, gm_n1225, gm_n158, in_19, gm_n2100, gm_n122);
	nand (gm_n2102, gm_n56, gm_n55, in_27, gm_n2101, gm_n182);
	nand (gm_n2103, gm_n2102, gm_n2099, gm_n2095);
	nor (gm_n2104, gm_n2082, gm_n2035, gm_n2031, gm_n2103, gm_n2092);
	nor (gm_n2105, gm_n669, gm_n62, gm_n61, gm_n670, gm_n284);
	nand (gm_n2106, gm_n121, gm_n158, gm_n58, gm_n2105, gm_n173);
	nor (gm_n2107, gm_n1112, gm_n55, in_27, gm_n2106, gm_n437);
	and (gm_n2108, gm_n199, gm_n65, gm_n62, gm_n883, gm_n174);
	nand (gm_n2109, gm_n459, in_23, gm_n58, gm_n2108, gm_n513);
	nor (gm_n2110, gm_n675, in_31, in_27, gm_n2109);
	nand (gm_n2111, gm_n110, gm_n63, gm_n124, gm_n402, gm_n144);
	nor (gm_n2112, gm_n188, gm_n76, gm_n73, gm_n2111, gm_n522);
	nand (gm_n2113, gm_n339, in_28, gm_n82, gm_n2112, gm_n263);
	nor (gm_n2114, gm_n2113, gm_n195);
	nor (gm_n2115, gm_n2114, gm_n2110, gm_n2107);
	nor (gm_n2116, gm_n599, in_12, in_8, gm_n1855, gm_n188);
	nand (gm_n2117, gm_n217, gm_n76, in_16, gm_n2116, gm_n477);
	nor (gm_n2118, gm_n195, in_28, in_24, gm_n2117, gm_n774);
	or (gm_n2119, gm_n116, gm_n63, in_8, gm_n282, gm_n178);
	nor (gm_n2120, gm_n249, in_20, in_16, gm_n2119, gm_n108);
	nand (gm_n2121, gm_n84, in_28, gm_n82, gm_n2120, gm_n263);
	nor (gm_n2122, gm_n2121, gm_n226);
	nor (gm_n2123, gm_n623, in_15, in_11, gm_n758, gm_n664);
	nand (gm_n2124, gm_n316, gm_n158, gm_n58, gm_n2123, gm_n455);
	nor (gm_n2125, gm_n1112, in_31, gm_n54, gm_n2124, gm_n423);
	nor (gm_n2126, gm_n2125, gm_n2122, gm_n2118);
	nand (gm_n2127, gm_n2104, gm_n2028, gm_n2025, gm_n2126, gm_n2115);
	nor (gm_n2128, gm_n664, gm_n753, gm_n447);
	nand (gm_n2129, gm_n123, in_15, gm_n61, gm_n2128, gm_n359);
	nor (gm_n2130, gm_n1225, gm_n158, gm_n58, gm_n2129, gm_n1112);
	nand (gm_n2131, gm_n308, gm_n55, in_27, gm_n2130);
	nor (gm_n2132, gm_n447, in_12, gm_n124, gm_n571, gm_n599);
	nand (gm_n2133, gm_n150, in_20, in_16, gm_n2132, gm_n521);
	nor (gm_n2134, gm_n224, in_28, gm_n82, gm_n2133, gm_n206);
	nand (gm_n2135, gm_n2134, gm_n81);
	nor (gm_n2136, gm_n151, gm_n115, gm_n70, gm_n469, gm_n124);
	and (gm_n2137, gm_n142, in_16, gm_n63, gm_n2136, gm_n242);
	and (gm_n2138, gm_n88, in_24, gm_n76, gm_n2137, gm_n235);
	nand (gm_n2139, gm_n225, gm_n84, gm_n83, gm_n2138);
	nand (gm_n2140, gm_n2139, gm_n2135, gm_n2131);
	nand (gm_n2141, gm_n112, in_1, gm_n94, in_4, gm_n68);
	nor (gm_n2142, gm_n345, gm_n2141);
	nand (gm_n2143, gm_n394, in_15, in_11, gm_n2142, gm_n1226);
	nor (gm_n2144, gm_n131, gm_n158, gm_n58, gm_n2143, gm_n393);
	nand (gm_n2145, gm_n182, in_31, in_27, gm_n2144, gm_n674);
	or (gm_n2146, gm_n553, in_16, in_12, gm_n1634, gm_n282);
	nor (gm_n2147, gm_n206, in_24, in_20, gm_n2146, gm_n476);
	nand (gm_n2148, gm_n367, gm_n81, in_28, gm_n2147);
	nand (gm_n2149, gm_n126, gm_n71, in_11, gm_n502);
	or (gm_n2150, gm_n303, gm_n58, gm_n62, gm_n2149, gm_n398);
	nor (gm_n2151, gm_n583, in_27, gm_n158, gm_n2150, gm_n514);
	nand (gm_n2152, gm_n2151, gm_n308, in_31);
	nand (gm_n2153, gm_n2152, gm_n2148, gm_n2145);
	nor (gm_n2154, gm_n2127, gm_n2021, gm_n2018, gm_n2153, gm_n2140);
	and (gm_n2155, gm_n207, in_12, gm_n124, gm_n1506, gm_n242);
	nand (gm_n2156, gm_n103, gm_n76, gm_n73, gm_n2155, gm_n521);
	nor (gm_n2157, gm_n140, gm_n83, gm_n82, gm_n2156, gm_n226);
	nand (gm_n2158, gm_n310, gm_n265, in_8);
	nor (gm_n2159, gm_n236, in_16, in_12, gm_n2158, gm_n599);
	nand (gm_n2160, gm_n107, gm_n82, in_20, gm_n2159, gm_n192);
	nor (gm_n2161, gm_n262, gm_n234, in_28, gm_n2160);
	and (gm_n2162, gm_n153, gm_n71, in_8, gm_n594);
	and (gm_n2163, gm_n121, in_19, gm_n62, gm_n2162, gm_n313);
	nand (gm_n2164, gm_n173, gm_n54, gm_n158, gm_n2163, gm_n309);
	nor (gm_n2165, gm_n2164, gm_n437, in_31);
	nor (gm_n2166, gm_n2165, gm_n2161, gm_n2157);
	nor (gm_n2167, gm_n109, in_16, in_12, gm_n776, gm_n154);
	nand (gm_n2168, gm_n88, gm_n82, gm_n76, gm_n2167, gm_n164);
	nor (gm_n2169, gm_n479, gm_n262, gm_n83, gm_n2168);
	nand (gm_n2170, gm_n703, gm_n218, gm_n124);
	nor (gm_n2171, gm_n374, gm_n73, in_12, gm_n2170, gm_n352);
	nand (gm_n2172, gm_n263, gm_n82, in_20, gm_n2171, gm_n521);
	nor (gm_n2173, gm_n248, gm_n234, gm_n83, gm_n2172);
	nor (gm_n2174, gm_n553, gm_n73, in_12, gm_n375, gm_n599);
	nand (gm_n2175, gm_n205, in_24, gm_n76, gm_n2174, gm_n477);
	nor (gm_n2176, gm_n684, gm_n774, gm_n83, gm_n2175);
	nor (gm_n2177, gm_n2176, gm_n2173, gm_n2169);
	nand (gm_n2178, gm_n2154, gm_n2015, gm_n2011, gm_n2177, gm_n2166);
	or (gm_n2179, gm_n249, in_16, in_12, gm_n266, gm_n282);
	nor (gm_n2180, gm_n104, gm_n82, in_20, gm_n2179, gm_n108);
	nand (gm_n2181, gm_n186, gm_n137, gm_n83, gm_n2180);
	not (gm_n2182, gm_n1180);
	nor (gm_n2183, in_9, gm_n124, gm_n151, gm_n535);
	nor (gm_n2184, in_12, gm_n61, in_10);
	nand (gm_n2185, gm_n404, gm_n105, in_13, gm_n2184, gm_n2183);
	nor (gm_n2186, gm_n2182, gm_n133, in_21, gm_n2185, gm_n1561);
	nand (gm_n2187, gm_n55, gm_n100, in_29, gm_n2186, gm_n408);
	nand (gm_n2188, gm_n208, gm_n127, gm_n124);
	or (gm_n2189, gm_n143, gm_n73, in_12, gm_n2188, gm_n288);
	nor (gm_n2190, gm_n520, in_24, in_20, gm_n2189, gm_n412);
	nand (gm_n2191, gm_n84, gm_n81, in_28, gm_n2190);
	nand (gm_n2192, gm_n2191, gm_n2187, gm_n2181);
	nand (gm_n2193, gm_n144, gm_n63, in_8, gm_n219, gm_n167);
	nor (gm_n2194, gm_n108, in_20, gm_n73, gm_n2193, gm_n109);
	nand (gm_n2195, gm_n139, gm_n83, in_24, gm_n2194, gm_n263);
	nor (gm_n2196, gm_n2195, gm_n185);
	nor (out_8, gm_n2192, gm_n2178, gm_n2006, gm_n2196);
	and (gm_n2198, gm_n199, in_12, in_8, gm_n588, gm_n264);
	and (gm_n2199, gm_n404, in_17, gm_n175, gm_n2198, gm_n1560);
	nand (gm_n2200, gm_n328, in_25, in_21, gm_n2199, gm_n539);
	nor (gm_n2201, gm_n55, gm_n100, gm_n80, gm_n2200);
	nand (gm_n2202, gm_n166, in_16, gm_n63, gm_n2136, gm_n256);
	nor (gm_n2203, gm_n108, gm_n82, gm_n76, gm_n2202, gm_n520);
	nand (gm_n2204, gm_n496, gm_n84, gm_n83, gm_n2203);
	and (gm_n2205, gm_n588, gm_n264, gm_n124);
	nand (gm_n2206, gm_n200, gm_n73, in_12, gm_n2205, gm_n340);
	nor (gm_n2207, gm_n108, in_24, in_20, gm_n2206, gm_n801);
	nand (gm_n2208, gm_n186, gm_n101, in_28, gm_n2207);
	not (gm_n2209, gm_n735);
	nor (gm_n2210, gm_n536, gm_n105, in_13, gm_n1126, gm_n767);
	nand (gm_n2211, gm_n651, gm_n133, in_21, gm_n2210, gm_n1560);
	nor (gm_n2212, gm_n55, gm_n100, gm_n80, gm_n2211, gm_n2209);
	and (gm_n2213, gm_n199, gm_n73, in_12, gm_n1887, gm_n446);
	nand (gm_n2214, gm_n141, gm_n82, in_20, gm_n2213, gm_n263);
	nor (gm_n2215, gm_n774, gm_n138, in_28, gm_n2214);
	nor (gm_n2216, gm_n152, gm_n63, gm_n124, gm_n2141, gm_n92);
	nand (gm_n2217, gm_n141, in_20, gm_n73, gm_n2216, gm_n446);
	nor (gm_n2218, gm_n140, gm_n83, in_24, gm_n2217, gm_n801);
	nand (gm_n2219, gm_n2218, gm_n496);
	or (gm_n2220, gm_n64, gm_n175, gm_n63, gm_n1387, gm_n154);
	or (gm_n2221, in_17, gm_n73, in_15, gm_n2220, in_18);
	nand (gm_n2222, in_21, gm_n76, gm_n58);
	nor (gm_n2223, gm_n640, in_26, in_22, gm_n2222, gm_n2221);
	nor (gm_n2224, in_29, gm_n83, gm_n54);
	nand (gm_n2225, gm_n2223, in_31, gm_n100, gm_n2224);
	nor (gm_n2226, gm_n571, gm_n152);
	and (gm_n2227, gm_n123, gm_n62, gm_n61, gm_n2226, gm_n930);
	nand (gm_n2228, gm_n121, in_23, gm_n58, gm_n2227, gm_n296);
	nor (gm_n2229, gm_n1112, gm_n55, gm_n54, gm_n2228, gm_n423);
	nor (gm_n2230, gm_n322, in_15, in_11, gm_n1201, gm_n398);
	nand (gm_n2231, gm_n334, gm_n158, in_19, gm_n2230, gm_n1042);
	nor (gm_n2232, gm_n1200, in_31, in_27, gm_n2231, gm_n838);
	or (gm_n2233, gm_n177, gm_n73, in_12, gm_n1117, gm_n282);
	nor (gm_n2234, gm_n89, gm_n82, gm_n76, gm_n2233, gm_n463);
	nand (gm_n2235, gm_n139, gm_n81, in_28, gm_n2234);
	nand (gm_n2236, gm_n153, gm_n63, in_8, gm_n973, gm_n176);
	nor (gm_n2237, gm_n165, in_20, in_16, gm_n2236, gm_n801);
	nand (gm_n2238, gm_n102, in_28, in_24, gm_n2237, gm_n213);
	and (gm_n2239, gm_n199, in_16, in_12, gm_n1499, gm_n166);
	nand (gm_n2240, gm_n90, in_24, gm_n76, gm_n2239, gm_n192);
	nor (gm_n2241, gm_n774, gm_n234, gm_n83, gm_n2240);
	and (gm_n2242, gm_n166, in_16, gm_n63, gm_n562, gm_n228);
	nand (gm_n2243, gm_n205, gm_n82, in_20, gm_n2242, gm_n270);
	nor (gm_n2244, gm_n248, gm_n234, in_28, gm_n2243);
	nand (gm_n2245, gm_n257, gm_n144, in_8);
	nor (gm_n2246, gm_n111, gm_n249, gm_n63, gm_n2245, gm_n613);
	nand (gm_n2247, gm_n296, in_23, gm_n58, gm_n2246, gm_n309);
	nor (gm_n2248, gm_n423, in_31, gm_n54, gm_n2247);
	nor (gm_n2249, gm_n360, gm_n62, gm_n61, gm_n1618, gm_n425);
	nand (gm_n2250, gm_n60, gm_n158, in_19, gm_n2249, gm_n296);
	nor (gm_n2251, gm_n57, in_31, gm_n54, gm_n2250);
	nor (gm_n2252, gm_n111, gm_n63, gm_n124, gm_n1527, gm_n374);
	nand (gm_n2253, gm_n90, gm_n76, gm_n73, gm_n2252, gm_n255);
	nor (gm_n2254, gm_n224, gm_n83, gm_n82, gm_n2253, gm_n684);
	nor (gm_n2255, gm_n2248, gm_n2244, gm_n2241, gm_n2254, gm_n2251);
	nand (gm_n2256, gm_n127, gm_n797, in_11, gm_n128);
	nor (gm_n2257, gm_n456, in_19, gm_n62, gm_n2256, gm_n623);
	nand (gm_n2258, gm_n358, in_27, gm_n158, gm_n2257, gm_n657);
	nor (gm_n2259, gm_n2258, gm_n357, gm_n55);
	nor (gm_n2260, gm_n360, gm_n58, gm_n62, gm_n996, gm_n425);
	nand (gm_n2261, gm_n309, in_27, in_23, gm_n2260, gm_n358);
	nor (gm_n2262, gm_n2261, gm_n612, gm_n55);
	nand (gm_n2263, gm_n243, gm_n144, in_8, gm_n426, gm_n256);
	nor (gm_n2264, gm_n796, in_19, gm_n62, gm_n2263, gm_n514);
	nand (gm_n2265, gm_n134, in_27, gm_n158, gm_n2264, gm_n306);
	nor (gm_n2266, gm_n2265, gm_n55);
	nor (gm_n2267, gm_n2266, gm_n2262, gm_n2259);
	nor (gm_n2268, gm_n796, in_15, in_11, gm_n1651, gm_n398);
	nand (gm_n2269, gm_n305, in_23, gm_n58, gm_n2268, gm_n316);
	nor (gm_n2270, gm_n357, gm_n55, gm_n54, gm_n2269);
	nor (gm_n2271, gm_n360, gm_n62, in_11, gm_n747, gm_n425);
	nand (gm_n2272, gm_n77, gm_n158, in_19, gm_n2271, gm_n134);
	nor (gm_n2273, gm_n618, in_31, in_27, gm_n2272);
	nand (gm_n2274, gm_n775, gm_n310);
	nor (gm_n2275, gm_n425, in_15, gm_n61, gm_n2274, gm_n664);
	nand (gm_n2276, gm_n174, in_23, gm_n58, gm_n2275, gm_n334);
	nor (gm_n2277, gm_n57, in_31, gm_n54, gm_n2276, gm_n1200);
	nor (gm_n2278, gm_n2277, gm_n2273, gm_n2270);
	nand (gm_n2279, gm_n2255, gm_n2238, gm_n2235, gm_n2278, gm_n2267);
	nand (gm_n2280, gm_n207, gm_n73, in_12, gm_n981, gm_n242);
	nor (gm_n2281, gm_n197, in_24, gm_n76, gm_n2280, gm_n801);
	nand (gm_n2282, gm_n225, gm_n186, gm_n83, gm_n2281);
	nand (gm_n2283, gm_n174, in_19, gm_n62, gm_n1999, gm_n1226);
	nor (gm_n2284, gm_n131, in_27, gm_n158, gm_n2283, gm_n977);
	nand (gm_n2285, gm_n2284, gm_n438, gm_n55);
	nand (gm_n2286, gm_n110, in_16, in_12, gm_n870, gm_n446);
	nor (gm_n2287, gm_n520, gm_n82, in_20, gm_n2286, gm_n463);
	nand (gm_n2288, gm_n139, gm_n81, in_28, gm_n2287);
	nand (gm_n2289, gm_n2288, gm_n2285, gm_n2282);
	or (gm_n2290, gm_n143, gm_n73, in_12, gm_n776, gm_n599);
	nor (gm_n2291, gm_n197, gm_n82, gm_n76, gm_n2290, gm_n630);
	nand (gm_n2292, gm_n339, gm_n81, in_28, gm_n2291);
	nand (gm_n2293, gm_n167, in_16, gm_n63, gm_n516, gm_n446);
	nor (gm_n2294, gm_n104, in_24, in_20, gm_n2293, gm_n463);
	nand (gm_n2295, gm_n496, gm_n102, in_28, gm_n2294);
	nand (gm_n2296, gm_n142, in_16, in_12, gm_n913, gm_n340);
	nor (gm_n2297, gm_n89, gm_n82, in_20, gm_n2296, gm_n197);
	nand (gm_n2298, gm_n213, gm_n139, in_28, gm_n2297);
	nand (gm_n2299, gm_n2298, gm_n2295, gm_n2292);
	nor (gm_n2300, gm_n2279, gm_n2232, gm_n2229, gm_n2299, gm_n2289);
	nor (gm_n2301, gm_n669, in_19, in_15, gm_n2149, gm_n393);
	nand (gm_n2302, gm_n296, gm_n54, gm_n158, gm_n2301, gm_n391);
	nor (gm_n2303, gm_n2302, gm_n357, in_31);
	nor (gm_n2304, gm_n584, gm_n62, gm_n61, gm_n664, gm_n623);
	nand (gm_n2305, gm_n121, gm_n158, in_19, gm_n2304, gm_n334);
	nor (gm_n2306, gm_n512, gm_n55, in_27, gm_n2305, gm_n357);
	nand (gm_n2307, gm_n515, gm_n208);
	nor (gm_n2308, gm_n111, gm_n63, gm_n124, gm_n2307, gm_n143);
	nand (gm_n2309, gm_n88, in_20, in_16, gm_n2308, gm_n477);
	nor (gm_n2310, gm_n214, gm_n83, gm_n82, gm_n2309, gm_n774);
	nor (gm_n2311, gm_n2310, gm_n2306, gm_n2303);
	nor (gm_n2312, gm_n109, gm_n73, in_12, gm_n1230, gm_n237);
	nand (gm_n2313, gm_n88, in_24, gm_n76, gm_n2312, gm_n270);
	nor (gm_n2314, gm_n479, gm_n774, in_28, gm_n2313);
	nor (gm_n2315, gm_n188, in_16, in_12, gm_n1019, gm_n352);
	nand (gm_n2316, gm_n107, in_24, gm_n76, gm_n2315, gm_n227);
	nor (gm_n2317, gm_n684, gm_n216, in_28, gm_n2316);
	nor (gm_n2318, gm_n236, in_16, gm_n63, gm_n1641, gm_n288);
	nand (gm_n2319, gm_n192, in_24, gm_n76, gm_n2318, gm_n521);
	nor (gm_n2320, gm_n684, gm_n224, gm_n83, gm_n2319);
	nor (gm_n2321, gm_n2320, gm_n2317, gm_n2314);
	nand (gm_n2322, gm_n2300, gm_n2225, gm_n2219, gm_n2321, gm_n2311);
	and (gm_n2323, gm_n594, gm_n310, in_11, gm_n730, gm_n622);
	nand (gm_n2324, gm_n359, gm_n58, in_15, gm_n2323, gm_n513);
	nor (gm_n2325, gm_n512, in_27, gm_n158, gm_n2324, gm_n612);
	nand (gm_n2326, gm_n2325, gm_n55);
	nand (gm_n2327, gm_n1137, gm_n264, gm_n124);
	or (gm_n2328, gm_n109, gm_n73, gm_n63, gm_n2327, gm_n154);
	nor (gm_n2329, gm_n187, in_24, gm_n76, gm_n2328, gm_n801);
	nand (gm_n2330, gm_n466, gm_n196, gm_n83, gm_n2329);
	nand (gm_n2331, gm_n200, gm_n73, gm_n63, gm_n784, gm_n340);
	nor (gm_n2332, gm_n104, in_24, gm_n76, gm_n2331, gm_n165);
	nand (gm_n2333, gm_n367, gm_n101, gm_n83, gm_n2332);
	nand (gm_n2334, gm_n2333, gm_n2330, gm_n2326);
	nor (gm_n2335, gm_n156, gm_n133, in_21, gm_n2009, gm_n532);
	nand (gm_n2336, gm_n55, gm_n100, gm_n80, gm_n2335, gm_n770);
	nand (gm_n2337, gm_n150, in_16, gm_n63, gm_n1173, gm_n242);
	nor (gm_n2338, gm_n108, in_24, gm_n76, gm_n2337, gm_n411);
	nand (gm_n2339, gm_n496, gm_n102, in_28, gm_n2338);
	nand (gm_n2340, gm_n207, in_16, gm_n63, gm_n709, gm_n256);
	nor (gm_n2341, gm_n187, in_24, in_20, gm_n2340, gm_n801);
	nand (gm_n2342, gm_n139, gm_n81, gm_n83, gm_n2341);
	nand (gm_n2343, gm_n2342, gm_n2339, gm_n2336);
	nor (gm_n2344, gm_n2322, gm_n2215, gm_n2212, gm_n2343, gm_n2334);
	nand (gm_n2345, gm_n588, gm_n218, in_8);
	nor (gm_n2346, gm_n249, in_16, gm_n63, gm_n2345, gm_n237);
	nand (gm_n2347, gm_n107, in_24, gm_n76, gm_n2346, gm_n227);
	nor (gm_n2348, gm_n216, gm_n214, gm_n83, gm_n2347);
	nand (gm_n2349, gm_n141, gm_n82, gm_n76, gm_n2137, gm_n255);
	nor (gm_n2350, gm_n214, gm_n85, gm_n83, gm_n2349);
	and (gm_n2351, gm_n123, gm_n62, in_11, gm_n1537, gm_n730);
	nand (gm_n2352, gm_n302, in_23, gm_n58, gm_n2351, gm_n358);
	nor (gm_n2353, gm_n1112, gm_n55, in_27, gm_n2352, gm_n612);
	nor (gm_n2354, gm_n2353, gm_n2350, gm_n2348);
	and (gm_n2355, gm_n107, in_20, gm_n73, gm_n1308, gm_n200);
	nand (gm_n2356, gm_n88, gm_n83, gm_n82, gm_n2355, gm_n466);
	nor (gm_n2357, gm_n2356, gm_n214);
	nor (gm_n2358, gm_n109, in_16, gm_n63, gm_n2032, gm_n599);
	nand (gm_n2359, gm_n88, gm_n82, in_20, gm_n2358, gm_n164);
	nor (gm_n2360, gm_n684, gm_n248, in_28, gm_n2359);
	nand (gm_n2361, in_6, in_5, in_4, gm_n320, in_7);
	nor (gm_n2362, gm_n623, gm_n62, gm_n61, gm_n2361, gm_n664);
	nand (gm_n2363, gm_n77, in_23, gm_n58, gm_n2362, gm_n302);
	nor (gm_n2364, gm_n57, in_31, in_27, gm_n2363, gm_n422);
	nor (gm_n2365, gm_n2364, gm_n2360, gm_n2357);
	nand (gm_n2366, gm_n2344, gm_n2208, gm_n2204, gm_n2365, gm_n2354);
	and (gm_n2367, gm_n228, in_12, in_8, gm_n594, gm_n264);
	nand (gm_n2368, gm_n107, in_20, in_16, gm_n2367, gm_n150);
	nor (gm_n2369, gm_n216, in_28, gm_n82, gm_n2368, gm_n630);
	nand (gm_n2370, gm_n2369, gm_n629);
	or (gm_n2371, gm_n432, in_15, in_11, gm_n1268, gm_n322);
	nor (gm_n2372, gm_n796, gm_n158, gm_n58, gm_n2371, gm_n335);
	nand (gm_n2373, gm_n182, in_31, in_27, gm_n2372, gm_n511);
	nand (gm_n2374, gm_n2022, in_15, in_11, gm_n730, gm_n622);
	nor (gm_n2375, gm_n452, gm_n158, in_19, gm_n2374, gm_n303);
	nand (gm_n2376, gm_n182, gm_n55, gm_n54, gm_n2375, gm_n337);
	nand (gm_n2377, gm_n2376, gm_n2373, gm_n2370);
	nand (gm_n2378, gm_n141, in_24, gm_n76, gm_n1571, gm_n227);
	nor (gm_n2379, gm_n368, gm_n185, in_28, gm_n2378);
	nor (out_9, gm_n2377, gm_n2366, gm_n2201, gm_n2379);
	nand (gm_n2381, gm_n394, gm_n311, gm_n127);
	nor (gm_n2382, gm_n303, gm_n62, in_11, gm_n2381, gm_n314);
	nand (gm_n2383, gm_n130, in_23, in_19, gm_n2382, gm_n657);
	nor (gm_n2384, gm_n675, gm_n55, gm_n54, gm_n2383);
	or (gm_n2385, gm_n143, gm_n63, in_8, gm_n384, gm_n288);
	nor (gm_n2386, gm_n411, gm_n76, gm_n73, gm_n2385, gm_n476);
	nand (gm_n2387, gm_n81, in_28, gm_n82, gm_n2386, gm_n215);
	nand (gm_n2388, gm_n310, gm_n228, gm_n124, gm_n620);
	or (gm_n2389, gm_n122, in_19, in_15, gm_n2388, gm_n363);
	nor (gm_n2390, gm_n431, gm_n54, in_23, gm_n2389, gm_n977);
	nand (gm_n2391, gm_n2390, gm_n306, in_31);
	nor (gm_n2392, gm_n143, in_20, gm_n73, gm_n1088, gm_n165);
	nand (gm_n2393, gm_n192, in_28, in_24, gm_n2392, gm_n466);
	nor (gm_n2394, gm_n2393, gm_n195);
	and (gm_n2395, gm_n110, gm_n73, gm_n63, gm_n879, gm_n207);
	nand (gm_n2396, gm_n141, gm_n82, gm_n76, gm_n2395, gm_n192);
	nor (gm_n2397, gm_n262, gm_n226, in_28, gm_n2396);
	nand (gm_n2398, gm_n176, gm_n73, in_12, gm_n448, gm_n340);
	nor (gm_n2399, gm_n187, in_24, in_20, gm_n2398, gm_n411);
	nand (gm_n2400, gm_n137, gm_n84, in_28, gm_n2399);
	nor (gm_n2401, in_7, gm_n115, gm_n70, gm_n469, gm_n124);
	nand (gm_n2402, gm_n199, in_16, in_12, gm_n2401, gm_n200);
	nor (gm_n2403, gm_n520, gm_n82, gm_n76, gm_n2402, gm_n412);
	nand (gm_n2404, gm_n496, gm_n466, in_28, gm_n2403);
	nor (gm_n2405, gm_n599, gm_n73, in_12, gm_n909, gm_n188);
	nand (gm_n2406, gm_n107, in_24, gm_n76, gm_n2405, gm_n263);
	nor (gm_n2407, gm_n684, gm_n248, in_28, gm_n2406);
	nand (gm_n2408, gm_n74, gm_n158, in_19, gm_n655, gm_n173);
	nor (gm_n2409, gm_n183, gm_n55, gm_n54, gm_n2408, gm_n838);
	or (gm_n2410, gm_n669, gm_n62, in_11, gm_n1479, gm_n395);
	nor (gm_n2411, gm_n514, gm_n158, gm_n58, gm_n2410, gm_n613);
	nand (gm_n2412, gm_n182, in_31, in_27, gm_n2411, gm_n511);
	nand (gm_n2413, gm_n446, in_16, in_12, gm_n1887, gm_n242);
	nor (gm_n2414, gm_n206, in_24, gm_n76, gm_n2413, gm_n463);
	nand (gm_n2415, gm_n339, gm_n137, in_28, gm_n2414);
	and (gm_n2416, gm_n340, gm_n74, gm_n62, gm_n516, gm_n698);
	nand (gm_n2417, gm_n513, gm_n158, gm_n58, gm_n2416, gm_n657);
	nor (gm_n2418, gm_n437, in_31, in_27, gm_n2417);
	nor (gm_n2419, gm_n322, in_15, in_11, gm_n1322, gm_n363);
	nand (gm_n2420, gm_n74, in_23, in_19, gm_n2419, gm_n358);
	nor (gm_n2421, gm_n437, in_31, in_27, gm_n2420, gm_n458);
	and (gm_n2422, gm_n142, in_12, in_8, gm_n1133, gm_n153);
	nand (gm_n2423, gm_n103, in_20, gm_n73, gm_n2422, gm_n164);
	nor (gm_n2424, gm_n216, gm_n83, in_24, gm_n2423, gm_n226);
	nor (gm_n2425, gm_n109, gm_n73, gm_n63, gm_n2170, gm_n288);
	nand (gm_n2426, gm_n192, gm_n82, gm_n76, gm_n2425, gm_n235);
	nor (gm_n2427, gm_n479, gm_n224, in_28, gm_n2426);
	and (gm_n2428, gm_n313, gm_n62, gm_n61, gm_n699, gm_n424);
	nand (gm_n2429, gm_n77, in_23, gm_n58, gm_n2428, gm_n392);
	nor (gm_n2430, gm_n512, gm_n55, in_27, gm_n2429, gm_n357);
	nor (gm_n2431, gm_n2424, gm_n2421, gm_n2418, gm_n2430, gm_n2427);
	and (gm_n2432, gm_n797, gm_n62, gm_n61, gm_n1626, gm_n698);
	nand (gm_n2433, gm_n130, gm_n158, gm_n58, gm_n2432, gm_n392);
	nor (gm_n2434, gm_n612, in_31, in_27, gm_n2433, gm_n977);
	nor (gm_n2435, gm_n670, gm_n62, gm_n61, gm_n2074, gm_n623);
	nand (gm_n2436, gm_n316, gm_n158, gm_n58, gm_n2435, gm_n1042);
	nor (gm_n2437, gm_n977, gm_n55, gm_n54, gm_n2436, gm_n675);
	and (gm_n2438, gm_n150, in_16, gm_n63, gm_n2012, gm_n167);
	nand (gm_n2439, gm_n164, in_24, in_20, gm_n2438, gm_n255);
	nor (gm_n2440, gm_n140, gm_n138, in_28, gm_n2439);
	nor (gm_n2441, gm_n2440, gm_n2437, gm_n2434);
	nor (gm_n2442, gm_n105, gm_n73, gm_n62, gm_n2220, gm_n106);
	nor (gm_n2443, gm_n86, gm_n76, in_19);
	nor (gm_n2444, in_25, gm_n82, gm_n158);
	nand (gm_n2445, gm_n2442, in_26, gm_n87, gm_n2444, gm_n2443);
	or (gm_n2446, in_29, in_28, in_27);
	nor (gm_n2447, gm_n2445, gm_n55, in_30, gm_n2446);
	nor (gm_n2448, gm_n599, gm_n73, gm_n63, gm_n1046, gm_n177);
	nand (gm_n2449, gm_n227, in_24, gm_n76, gm_n2448, gm_n235);
	nor (gm_n2450, gm_n248, gm_n138, gm_n83, gm_n2449);
	nand (gm_n2451, gm_n128, gm_n189, in_11, gm_n698, gm_n930);
	nor (gm_n2452, gm_n122, gm_n58, in_15, gm_n2451, gm_n317);
	nand (gm_n2453, gm_n390, gm_n54, in_23, gm_n2452, gm_n391);
	nor (gm_n2454, gm_n2453, in_31);
	nor (gm_n2455, gm_n2454, gm_n2450, gm_n2447);
	nand (gm_n2456, gm_n2431, gm_n2415, gm_n2412, gm_n2455, gm_n2441);
	and (gm_n2457, gm_n110, in_12, in_8, gm_n310, gm_n257);
	nand (gm_n2458, gm_n91, gm_n76, in_16, gm_n2457, gm_n235);
	nor (gm_n2459, gm_n104, gm_n83, gm_n82, gm_n2458, gm_n774);
	nand (gm_n2460, gm_n2459, gm_n137);
	or (gm_n2461, gm_n188, in_16, in_12, gm_n1405, gm_n288);
	nor (gm_n2462, gm_n566, gm_n82, in_20, gm_n2461, gm_n522);
	nand (gm_n2463, gm_n139, gm_n101, in_28, gm_n2462);
	nor (gm_n2464, gm_n105, in_16, gm_n62);
	nand (gm_n2465, gm_n484, in_14, gm_n61, gm_n2464, gm_n485);
	nor (gm_n2466, gm_n490, gm_n87, gm_n106, gm_n2465, gm_n638);
	nand (gm_n2467, in_31, gm_n100, gm_n59, gm_n2466, gm_n1897);
	nand (gm_n2468, gm_n2467, gm_n2463, gm_n2460);
	nand (gm_n2469, gm_n207, gm_n73, in_12, gm_n866, gm_n340);
	nor (gm_n2470, gm_n520, gm_n82, gm_n76, gm_n2469, gm_n412);
	nand (gm_n2471, gm_n215, gm_n81, in_28, gm_n2470);
	nand (gm_n2472, gm_n164, gm_n76, gm_n73, gm_n2367, gm_n446);
	nor (gm_n2473, gm_n224, in_28, gm_n82, gm_n2472, gm_n566);
	nand (gm_n2474, gm_n2473, gm_n81);
	nand (gm_n2475, gm_n91, gm_n73, gm_n63, gm_n866, gm_n228);
	nor (gm_n2476, gm_n566, gm_n82, gm_n76, gm_n2475, gm_n463);
	nand (gm_n2477, gm_n139, gm_n101, gm_n83, gm_n2476);
	nand (gm_n2478, gm_n2477, gm_n2474, gm_n2471);
	nor (gm_n2479, gm_n2456, gm_n2409, gm_n2407, gm_n2478, gm_n2468);
	nor (gm_n2480, gm_n92, in_16, gm_n63, gm_n2158, gm_n374);
	nand (gm_n2481, gm_n235, gm_n82, gm_n76, gm_n2480, gm_n263);
	nor (gm_n2482, gm_n479, gm_n224, gm_n83, gm_n2481);
	nor (gm_n2483, gm_n374, gm_n73, in_12, gm_n1405, gm_n282);
	nand (gm_n2484, gm_n90, gm_n82, in_20, gm_n2483, gm_n263);
	nor (gm_n2485, gm_n368, gm_n214, gm_n83, gm_n2484);
	and (gm_n2486, gm_n731, gm_n310, in_8);
	and (gm_n2487, gm_n167, gm_n73, gm_n63, gm_n2486, gm_n176);
	nand (gm_n2488, gm_n141, gm_n82, in_20, gm_n2487, gm_n205);
	nor (gm_n2489, gm_n684, gm_n140, gm_n83, gm_n2488);
	nor (gm_n2490, gm_n2489, gm_n2485, gm_n2482);
	nand (gm_n2491, gm_n145, in_4, gm_n68, gm_n310);
	nor (gm_n2492, gm_n669, in_15, gm_n61, gm_n2491, gm_n322);
	nand (gm_n2493, gm_n74, gm_n158, gm_n58, gm_n2492, gm_n130);
	nor (gm_n2494, gm_n618, gm_n55, gm_n54, gm_n2493, gm_n422);
	nor (gm_n2495, gm_n599, gm_n73, in_12, gm_n2188, gm_n177);
	nand (gm_n2496, gm_n141, gm_n82, gm_n76, gm_n2495, gm_n205);
	nor (gm_n2497, gm_n195, gm_n85, in_28, gm_n2496);
	and (gm_n2498, gm_n169, in_16, gm_n63, gm_n256, gm_n207);
	nand (gm_n2499, gm_n141, in_24, gm_n76, gm_n2498, gm_n205);
	nor (gm_n2500, gm_n684, gm_n248, in_28, gm_n2499);
	nor (gm_n2501, gm_n2500, gm_n2497, gm_n2494);
	nand (gm_n2502, gm_n2479, gm_n2404, gm_n2400, gm_n2501, gm_n2490);
	nand (gm_n2503, gm_n446, in_16, gm_n63, gm_n346, gm_n256);
	nor (gm_n2504, gm_n187, in_24, in_20, gm_n2503, gm_n206);
	nand (gm_n2505, gm_n213, gm_n186, in_28, gm_n2504);
	or (gm_n2506, gm_n92, in_15, in_8, gm_n1034, gm_n314);
	nor (gm_n2507, gm_n331, gm_n158, gm_n58, gm_n2506, gm_n335);
	nand (gm_n2508, gm_n60, gm_n55, gm_n54, gm_n2507, gm_n438);
	and (gm_n2509, gm_n127, gm_n63, gm_n124, gm_n731, gm_n228);
	nand (gm_n2510, gm_n91, in_20, in_16, gm_n2509, gm_n521);
	nor (gm_n2511, gm_n566, in_28, gm_n82, gm_n2510, gm_n262);
	nand (gm_n2512, gm_n2511, gm_n496);
	nand (gm_n2513, gm_n2512, gm_n2508, gm_n2505);
	and (gm_n2514, in_7, gm_n115, in_5, gm_n361, gm_n124);
	nand (gm_n2515, gm_n91, gm_n73, gm_n63, gm_n2514, gm_n228);
	nor (gm_n2516, gm_n104, gm_n82, gm_n76, gm_n2515, gm_n463);
	nand (gm_n2517, gm_n466, gm_n213, gm_n83, gm_n2516);
	nand (gm_n2518, gm_n200, gm_n76, gm_n73, gm_n1300, gm_n270);
	nor (gm_n2519, gm_n89, gm_n83, in_24, gm_n2518, gm_n140);
	nand (gm_n2520, gm_n2519, gm_n225);
	and (gm_n2521, gm_n127, gm_n63, gm_n124, gm_n289, gm_n167);
	nand (gm_n2522, gm_n200, gm_n76, in_16, gm_n2521, gm_n164);
	nor (gm_n2523, gm_n224, in_28, gm_n82, gm_n2522, gm_n801);
	nand (gm_n2524, gm_n2523, gm_n101);
	nand (gm_n2525, gm_n2524, gm_n2520, gm_n2517);
	nor (gm_n2526, gm_n2502, gm_n2397, gm_n2394, gm_n2525, gm_n2513);
	and (gm_n2527, gm_n107, gm_n76, gm_n73, gm_n2132, gm_n176);
	nand (gm_n2528, gm_n217, in_28, in_24, gm_n2527, gm_n466);
	nor (gm_n2529, gm_n2528, gm_n185);
	nor (gm_n2530, gm_n725, gm_n62, gm_n61, gm_n991, gm_n758);
	nand (gm_n2531, gm_n334, gm_n158, gm_n58, gm_n2530, gm_n359);
	nor (gm_n2532, gm_n57, in_31, gm_n54, gm_n2531, gm_n512);
	and (gm_n2533, gm_n91, in_16, gm_n63, gm_n1350, gm_n110);
	nand (gm_n2534, gm_n255, in_24, gm_n76, gm_n2533, gm_n477);
	nor (gm_n2535, gm_n195, gm_n140, gm_n83, gm_n2534);
	nor (gm_n2536, gm_n2535, gm_n2532, gm_n2529);
	and (gm_n2537, gm_n123, in_15, gm_n61, gm_n1081, gm_n394);
	nand (gm_n2538, gm_n173, gm_n158, gm_n58, gm_n2537, gm_n455);
	nor (gm_n2539, gm_n57, gm_n55, gm_n54, gm_n2538, gm_n183);
	and (gm_n2540, gm_n123, gm_n62, in_11, gm_n1760, gm_n930);
	nand (gm_n2541, gm_n334, gm_n158, in_19, gm_n2540, gm_n1042);
	nor (gm_n2542, gm_n57, gm_n55, in_27, gm_n2541, gm_n512);
	nand (gm_n2543, gm_n1137, gm_n310, gm_n124);
	nor (gm_n2544, gm_n109, in_16, in_12, gm_n2543, gm_n282);
	nand (gm_n2545, gm_n90, in_24, in_20, gm_n2544, gm_n263);
	nor (gm_n2546, gm_n248, gm_n138, gm_n83, gm_n2545);
	nor (gm_n2547, gm_n2546, gm_n2542, gm_n2539);
	nand (gm_n2548, gm_n2526, gm_n2391, gm_n2387, gm_n2547, gm_n2536);
	or (gm_n2549, gm_n669, in_19, in_15, gm_n614, gm_n393);
	nor (gm_n2550, gm_n458, gm_n54, in_23, gm_n2549, gm_n514);
	nand (gm_n2551, gm_n2550, gm_n438, in_31);
	or (gm_n2552, gm_n288, in_15, gm_n124, gm_n1527, gm_n363);
	nor (gm_n2553, gm_n452, in_23, in_19, gm_n2552, gm_n303);
	nand (gm_n2554, gm_n182, in_31, gm_n54, gm_n2553, gm_n308);
	nor (gm_n2555, gm_n971, gm_n178, gm_n124);
	nand (gm_n2556, gm_n166, gm_n73, gm_n63, gm_n2555, gm_n340);
	nor (gm_n2557, gm_n630, in_24, gm_n76, gm_n2556, gm_n522);
	nand (gm_n2558, gm_n225, gm_n102, gm_n83, gm_n2557);
	nand (gm_n2559, gm_n2558, gm_n2554, gm_n2551);
	and (gm_n2560, gm_n123, gm_n62, in_11, gm_n1545, gm_n1042);
	nand (gm_n2561, gm_n173, gm_n158, gm_n58, gm_n2560, gm_n459);
	nor (gm_n2562, gm_n357, in_31, in_27, gm_n2561);
	nor (out_10, gm_n2559, gm_n2548, gm_n2384, gm_n2562);
	nor (gm_n2564, gm_n154, in_12, in_8, gm_n1805, gm_n188);
	nand (gm_n2565, gm_n141, gm_n76, in_16, gm_n2564, gm_n263);
	nor (gm_n2566, gm_n214, gm_n83, gm_n82, gm_n2565, gm_n368);
	nor (gm_n2567, gm_n383, gm_n972, gm_n124);
	nand (gm_n2568, gm_n199, gm_n73, gm_n63, gm_n2567, gm_n446);
	nor (gm_n2569, gm_n187, gm_n82, in_20, gm_n2568, gm_n520);
	nand (gm_n2570, gm_n339, gm_n137, gm_n83, gm_n2569);
	or (gm_n2571, gm_n314, in_19, in_15, gm_n2056, gm_n360);
	nor (gm_n2572, gm_n131, gm_n54, gm_n158, gm_n2571, gm_n583);
	nand (gm_n2573, gm_n2572, gm_n511, gm_n55);
	nor (gm_n2574, gm_n143, gm_n73, in_12, gm_n1686, gm_n288);
	nand (gm_n2575, gm_n88, gm_n82, gm_n76, gm_n2574, gm_n90);
	nor (gm_n2576, gm_n226, gm_n140, in_28, gm_n2575);
	nor (gm_n2577, gm_n670, gm_n2141, gm_n447);
	and (gm_n2578, gm_n698, gm_n62, gm_n61, gm_n2577, gm_n455);
	nand (gm_n2579, gm_n296, gm_n158, in_19, gm_n2578, gm_n657);
	nor (gm_n2580, gm_n618, in_31, in_27, gm_n2579);
	nor (gm_n2581, gm_n151, gm_n115, gm_n70, gm_n114);
	nand (gm_n2582, gm_n698, gm_n62, gm_n61, gm_n2581, gm_n424);
	nor (gm_n2583, gm_n297, in_23, in_19, gm_n2582, gm_n456);
	nand (gm_n2584, gm_n459, in_31, in_27, gm_n2583, gm_n511);
	nor (gm_n2585, gm_n352, gm_n63, gm_n124, gm_n383, gm_n229);
	and (gm_n2586, gm_n1178, gm_n105, gm_n175, gm_n2585, gm_n1560);
	and (gm_n2587, gm_n328, gm_n133, gm_n86, gm_n2586, gm_n769);
	nand (gm_n2588, in_31, gm_n100, in_29, gm_n2587);
	or (gm_n2589, gm_n483, gm_n151);
	nor (gm_n2590, gm_n125, gm_n62, gm_n61, gm_n2589, gm_n398);
	nand (gm_n2591, gm_n334, in_23, in_19, gm_n2590, gm_n392);
	nor (gm_n2592, gm_n357, in_31, gm_n54, gm_n2591, gm_n422);
	nor (gm_n2593, gm_n599, gm_n73, gm_n63, gm_n2327, gm_n177);
	nand (gm_n2594, gm_n103, in_24, gm_n76, gm_n2593, gm_n107);
	nor (gm_n2595, gm_n216, gm_n214, gm_n83, gm_n2594);
	nand (gm_n2596, gm_n207, in_16, in_12, gm_n685, gm_n340);
	nor (gm_n2597, gm_n89, in_24, in_20, gm_n2596, gm_n165);
	nand (gm_n2598, gm_n466, gm_n213, gm_n83, gm_n2597);
	nor (gm_n2599, gm_n92, in_12, in_8, gm_n298, gm_n447);
	nand (gm_n2600, gm_n141, gm_n76, in_16, gm_n2599, gm_n142);
	nor (gm_n2601, gm_n104, gm_n83, in_24, gm_n2600, gm_n140);
	nand (gm_n2602, gm_n2601, gm_n81);
	nor (gm_n2603, gm_n432, gm_n62, in_11, gm_n671, gm_n725);
	nand (gm_n2604, gm_n173, gm_n158, gm_n58, gm_n2603, gm_n392);
	nor (gm_n2605, gm_n183, gm_n55, gm_n54, gm_n2604, gm_n437);
	nand (gm_n2606, gm_n358, in_23, gm_n58, gm_n1277, gm_n359);
	nor (gm_n2607, gm_n422, gm_n55, gm_n54, gm_n2606, gm_n437);
	nor (gm_n2608, gm_n249, gm_n73, in_12, gm_n2188, gm_n154);
	nand (gm_n2609, gm_n192, gm_n82, gm_n76, gm_n2608, gm_n477);
	nor (gm_n2610, gm_n479, gm_n85, gm_n83, gm_n2609);
	nor (gm_n2611, gm_n363, gm_n62, in_11, gm_n1272, gm_n664);
	nand (gm_n2612, gm_n130, gm_n158, gm_n58, gm_n2611, gm_n359);
	nor (gm_n2613, gm_n183, in_31, gm_n54, gm_n2612, gm_n612);
	nand (gm_n2614, gm_n256, in_12, in_8, gm_n594, gm_n264);
	nor (gm_n2615, gm_n553, in_20, gm_n73, gm_n2614, gm_n463);
	nand (gm_n2616, gm_n139, gm_n83, gm_n82, gm_n2615, gm_n192);
	nor (gm_n2617, gm_n2616, gm_n214);
	nor (gm_n2618, gm_n2610, gm_n2607, gm_n2605, gm_n2617, gm_n2613);
	nor (gm_n2619, gm_n177, gm_n73, in_12, gm_n1263, gm_n288);
	nand (gm_n2620, gm_n235, gm_n82, gm_n76, gm_n2619, gm_n263);
	nor (gm_n2621, gm_n195, gm_n140, in_28, gm_n2620);
	nor (gm_n2622, gm_n92, gm_n73, in_12, gm_n1795, gm_n143);
	nand (gm_n2623, gm_n255, gm_n82, in_20, gm_n2622, gm_n270);
	nor (gm_n2624, gm_n774, gm_n214, gm_n83, gm_n2623);
	nor (gm_n2625, gm_n374, gm_n73, gm_n63, gm_n2345, gm_n282);
	nand (gm_n2626, gm_n88, in_24, in_20, gm_n2625, gm_n477);
	nor (gm_n2627, gm_n224, gm_n185, in_28, gm_n2626);
	nor (gm_n2628, gm_n2627, gm_n2624, gm_n2621);
	nor (gm_n2629, gm_n249, in_12, in_8, gm_n2307, gm_n92);
	nand (gm_n2630, gm_n103, in_20, gm_n73, gm_n2629, gm_n235);
	nor (gm_n2631, gm_n234, gm_n83, gm_n82, gm_n2630, gm_n216);
	nor (gm_n2632, gm_n599, gm_n73, gm_n63, gm_n1296, gm_n177);
	nand (gm_n2633, gm_n192, gm_n82, in_20, gm_n2632, gm_n235);
	nor (gm_n2634, gm_n195, gm_n140, gm_n83, gm_n2633);
	or (gm_n2635, gm_n111, in_12, gm_n124, gm_n447, gm_n114);
	nor (gm_n2636, gm_n187, in_20, in_16, gm_n2635, gm_n374);
	nand (gm_n2637, gm_n102, in_28, in_24, gm_n2636, gm_n103);
	nor (gm_n2638, gm_n2637, gm_n195);
	nor (gm_n2639, gm_n2638, gm_n2634, gm_n2631);
	nand (gm_n2640, gm_n2618, gm_n2602, gm_n2598, gm_n2639, gm_n2628);
	or (gm_n2641, gm_n249, gm_n73, gm_n63, gm_n353, gm_n288);
	nor (gm_n2642, gm_n187, in_24, gm_n76, gm_n2641, gm_n801);
	nand (gm_n2643, gm_n225, gm_n215, gm_n83, gm_n2642);
	nor (gm_n2644, gm_n111, gm_n63, in_8, gm_n971, gm_n168);
	nand (gm_n2645, gm_n200, gm_n76, gm_n73, gm_n2644, gm_n521);
	nor (gm_n2646, gm_n248, in_28, gm_n82, gm_n2645, gm_n411);
	nand (gm_n2647, gm_n2646, gm_n101);
	nand (gm_n2648, gm_n91, in_16, gm_n63, gm_n1994, gm_n228);
	nor (gm_n2649, gm_n197, in_24, in_20, gm_n2648, gm_n801);
	nand (gm_n2650, gm_n367, gm_n101, gm_n83, gm_n2649);
	nand (gm_n2651, gm_n2650, gm_n2647, gm_n2643);
	nor (gm_n2652, gm_n972, gm_n93);
	nand (gm_n2653, gm_n797, in_15, in_11, gm_n2652, gm_n931);
	nor (gm_n2654, gm_n431, in_23, gm_n58, gm_n2653, gm_n456);
	nand (gm_n2655, gm_n306, in_31, gm_n54, gm_n2654, gm_n459);
	nand (gm_n2656, gm_n995, in_15, in_11, gm_n2226, gm_n698);
	nor (gm_n2657, gm_n131, gm_n158, in_19, gm_n2656, gm_n303);
	nand (gm_n2658, gm_n305, in_31, gm_n54, gm_n2657, gm_n337);
	nand (gm_n2659, gm_n199, gm_n73, gm_n63, gm_n1055, gm_n166);
	nor (gm_n2660, gm_n411, in_24, in_20, gm_n2659, gm_n522);
	nand (gm_n2661, gm_n339, gm_n137, in_28, gm_n2660);
	nand (gm_n2662, gm_n2661, gm_n2658, gm_n2655);
	nor (gm_n2663, gm_n2640, gm_n2595, gm_n2592, gm_n2662, gm_n2651);
	nor (gm_n2664, gm_n177, gm_n73, gm_n63, gm_n1019, gm_n282);
	nand (gm_n2665, gm_n205, in_24, in_20, gm_n2664, gm_n270);
	nor (gm_n2666, gm_n214, gm_n248, in_28, gm_n2665);
	nand (gm_n2667, gm_n151, gm_n115, in_5, gm_n361, gm_n124);
	nor (gm_n2668, gm_n92, in_16, in_12, gm_n2667, gm_n143);
	nand (gm_n2669, gm_n88, in_24, gm_n76, gm_n2668, gm_n107);
	nor (gm_n2670, gm_n774, gm_n185, gm_n83, gm_n2669);
	nor (gm_n2671, gm_n92, in_16, gm_n63, gm_n952, gm_n553);
	nand (gm_n2672, gm_n103, gm_n82, in_20, gm_n2671, gm_n477);
	nor (gm_n2673, gm_n479, gm_n140, gm_n83, gm_n2672);
	nor (gm_n2674, gm_n2673, gm_n2670, gm_n2666);
	nor (gm_n2675, gm_n284, in_15, in_11, gm_n425, gm_n670);
	nand (gm_n2676, gm_n74, in_23, gm_n58, gm_n2675, gm_n173);
	nor (gm_n2677, gm_n357, gm_n55, in_27, gm_n2676, gm_n422);
	or (gm_n2678, gm_n433, gm_n93, gm_n61, gm_n548, gm_n425);
	nor (gm_n2679, gm_n131, gm_n58, gm_n62, gm_n2678, gm_n456);
	nand (gm_n2680, gm_n182, gm_n54, in_23, gm_n2679, gm_n306);
	nor (gm_n2681, gm_n2680, in_31);
	or (gm_n2682, gm_n971, gm_n229);
	nor (gm_n2683, gm_n322, in_15, in_11, gm_n2682, gm_n363);
	nand (gm_n2684, gm_n130, gm_n158, in_19, gm_n2683, gm_n455);
	nor (gm_n2685, gm_n1200, gm_n55, in_27, gm_n2684, gm_n437);
	nor (gm_n2686, gm_n2685, gm_n2681, gm_n2677);
	nand (gm_n2687, gm_n2663, gm_n2588, gm_n2584, gm_n2686, gm_n2674);
	or (gm_n2688, gm_n314, gm_n62, gm_n61, gm_n554, gm_n395);
	nor (gm_n2689, gm_n393, gm_n158, in_19, gm_n2688, gm_n514);
	nand (gm_n2690, gm_n56, in_31, in_27, gm_n2689, gm_n305);
	nor (gm_n2691, gm_n95, gm_n63, in_8, gm_n971, gm_n282);
	nand (gm_n2692, gm_n200, gm_n76, in_16, gm_n2691, gm_n235);
	nor (gm_n2693, gm_n248, in_28, in_24, gm_n2692, gm_n630);
	nand (gm_n2694, gm_n2693, gm_n629);
	nand (gm_n2695, gm_n123, in_15, in_11, gm_n1626, gm_n930);
	nor (gm_n2696, gm_n131, gm_n158, gm_n58, gm_n2695, gm_n331);
	nand (gm_n2697, gm_n182, gm_n55, gm_n54, gm_n2696, gm_n674);
	nand (gm_n2698, gm_n2697, gm_n2694, gm_n2690);
	nor (gm_n2699, gm_n971, in_12, in_8, gm_n548, gm_n288);
	nand (gm_n2700, gm_n141, gm_n76, gm_n73, gm_n2699, gm_n166);
	nor (gm_n2701, gm_n206, gm_n83, in_24, gm_n2700, gm_n774);
	nand (gm_n2702, gm_n2701, gm_n101);
	nand (gm_n2703, gm_n392, gm_n199, in_15, gm_n883, gm_n622);
	nor (gm_n2704, gm_n1112, in_23, in_19, gm_n2703, gm_n335);
	nand (gm_n2705, gm_n56, in_31, gm_n54, gm_n2704);
	nor (gm_n2706, gm_n229, gm_n63, in_8, gm_n345, gm_n237);
	nand (gm_n2707, gm_n107, gm_n76, gm_n73, gm_n2706, gm_n166);
	nor (gm_n2708, gm_n411, in_28, gm_n82, gm_n2707, gm_n368);
	nand (gm_n2709, gm_n2708, gm_n629);
	nand (gm_n2710, gm_n2709, gm_n2705, gm_n2702);
	nor (gm_n2711, gm_n2687, gm_n2580, gm_n2576, gm_n2710, gm_n2698);
	or (gm_n2712, gm_n237, in_12, in_8, gm_n548, gm_n971);
	nor (gm_n2713, gm_n553, gm_n76, gm_n73, gm_n2712, gm_n165);
	nand (gm_n2714, gm_n186, in_28, gm_n82, gm_n2713, gm_n192);
	nor (gm_n2715, gm_n2714, gm_n185);
	nor (gm_n2716, gm_n109, in_16, gm_n63, gm_n1100, gm_n599);
	nand (gm_n2717, gm_n103, gm_n82, in_20, gm_n2716, gm_n235);
	nor (gm_n2718, gm_n224, gm_n234, in_28, gm_n2717);
	and (gm_n2719, gm_n91, in_16, in_12, gm_n754, gm_n242);
	nand (gm_n2720, gm_n227, gm_n82, gm_n76, gm_n2719, gm_n477);
	nor (gm_n2721, gm_n226, gm_n216, in_28, gm_n2720);
	nor (gm_n2722, gm_n2721, gm_n2718, gm_n2715);
	nor (gm_n2723, in_16, in_15);
	and (gm_n2724, gm_n2723, in_14);
	and (gm_n2725, gm_n405, in_17, gm_n175, gm_n2724, gm_n2198);
	nand (gm_n2726, gm_n769, gm_n133, in_21, gm_n2725);
	nor (gm_n2727, in_31, in_30, gm_n80, gm_n2726, gm_n1050);
	and (gm_n2728, gm_n1840, gm_n105, in_13, gm_n2007, gm_n1558);
	and (gm_n2729, gm_n159, in_25, gm_n86, gm_n2728, gm_n325);
	and (gm_n2730, gm_n55, in_30, in_29, gm_n2729, gm_n328);
	nor (gm_n2731, gm_n125, in_15, gm_n61, gm_n1252, gm_n425);
	nand (gm_n2732, gm_n130, gm_n158, in_19, gm_n2731, gm_n455);
	nor (gm_n2733, gm_n512, in_31, gm_n54, gm_n2732, gm_n618);
	nor (gm_n2734, gm_n2733, gm_n2730, gm_n2727);
	nand (gm_n2735, gm_n2711, gm_n2573, gm_n2570, gm_n2734, gm_n2722);
	nand (gm_n2736, gm_n126, in_15, in_11, gm_n1760, gm_n698);
	nor (gm_n2737, gm_n452, gm_n158, gm_n58, gm_n2736, gm_n456);
	nand (gm_n2738, gm_n134, gm_n55, in_27, gm_n2737, gm_n390);
	or (gm_n2739, gm_n143, in_16, gm_n63, gm_n1234, gm_n352);
	nor (gm_n2740, gm_n89, in_24, in_20, gm_n2739, gm_n197);
	nand (gm_n2741, gm_n339, gm_n101, in_28, gm_n2740);
	or (gm_n2742, gm_n553, gm_n73, in_12, gm_n1634, gm_n288);
	nor (gm_n2743, gm_n187, in_24, gm_n76, gm_n2742, gm_n411);
	nand (gm_n2744, gm_n215, gm_n196, gm_n83, gm_n2743);
	nand (gm_n2745, gm_n2744, gm_n2741, gm_n2738);
	nor (gm_n2746, gm_n92, in_16, gm_n63, gm_n2170, gm_n553);
	nand (gm_n2747, gm_n88, in_24, in_20, gm_n2746, gm_n477);
	nor (gm_n2748, gm_n262, gm_n195, in_28, gm_n2747);
	nor (out_11, gm_n2745, gm_n2735, gm_n2566, gm_n2748);
	not (gm_n2750, t_3);
	nor (gm_n2751, gm_n154, gm_n73, gm_n63, gm_n1059, gm_n236);
	and (gm_n2752, gm_n103, in_24, gm_n76, gm_n2751, gm_n164);
	and (gm_n2753, gm_n367, gm_n81, in_28, gm_n2752);
	nand (gm_n2754, gm_n446, in_16, gm_n63, gm_n1245, gm_n340);
	nor (gm_n2755, gm_n630, in_24, gm_n76, gm_n2754, gm_n412);
	nand (gm_n2756, gm_n215, gm_n81, gm_n83, gm_n2755);
	nand (gm_n2757, gm_n110, in_16, in_12, gm_n1015, gm_n150);
	nor (gm_n2758, gm_n801, in_24, gm_n76, gm_n2757, gm_n476);
	nand (gm_n2759, gm_n339, gm_n101, gm_n83, gm_n2758);
	nor (gm_n2760, gm_n249, gm_n76, gm_n73, gm_n2712, gm_n522);
	nand (gm_n2761, gm_n84, gm_n83, gm_n82, gm_n2760, gm_n88);
	nor (gm_n2762, gm_n2761, gm_n684);
	nor (gm_n2763, gm_n314, in_15, in_11, gm_n554, gm_n322);
	nand (gm_n2764, gm_n296, gm_n158, in_19, gm_n2763, gm_n1042);
	nor (gm_n2765, gm_n512, gm_n55, gm_n54, gm_n2764, gm_n437);
	and (gm_n2766, gm_n394, gm_n128, gm_n189);
	nand (gm_n2767, gm_n302, gm_n62, gm_n61, gm_n2766, gm_n698);
	nor (gm_n2768, gm_n183, gm_n158, gm_n58, gm_n2767, gm_n335);
	nand (gm_n2769, gm_n511, gm_n55, gm_n54, gm_n2768);
	and (gm_n2770, gm_n126, in_15, in_11, gm_n2652, gm_n313);
	nand (gm_n2771, gm_n173, in_23, in_19, gm_n2770, gm_n455);
	or (gm_n2772, gm_n1112, in_31, in_27, gm_n2771, gm_n423);
	nor (gm_n2773, gm_n92, gm_n73, gm_n63, gm_n1634, gm_n553);
	nand (gm_n2774, gm_n103, in_24, gm_n76, gm_n2773, gm_n164);
	nor (gm_n2775, gm_n684, gm_n368, in_28, gm_n2774);
	nor (gm_n2776, gm_n725, in_15, in_11, gm_n1272, gm_n991);
	nand (gm_n2777, gm_n173, gm_n158, gm_n58, gm_n2776, gm_n359);
	nor (gm_n2778, gm_n612, in_31, in_27, gm_n2777, gm_n458);
	nor (gm_n2779, gm_n282, gm_n62, gm_n124, gm_n991, gm_n384);
	nand (gm_n2780, gm_n77, in_23, in_19, gm_n2779, gm_n455);
	or (gm_n2781, gm_n422, in_31, gm_n54, gm_n2780, gm_n675);
	nor (gm_n2782, gm_n154, gm_n73, in_12, gm_n1772, gm_n188);
	and (gm_n2783, gm_n107, gm_n82, gm_n76, gm_n2782, gm_n205);
	nand (gm_n2784, gm_n496, gm_n186, in_28, gm_n2783);
	and (gm_n2785, gm_n142, gm_n73, gm_n63, gm_n1142, gm_n228);
	nand (gm_n2786, gm_n141, in_24, gm_n76, gm_n2785, gm_n263);
	nor (gm_n2787, gm_n684, gm_n216, in_28, gm_n2786);
	or (gm_n2788, gm_n73, gm_n62, in_14, gm_n1606, in_17);
	or (gm_n2789, gm_n157, gm_n133, gm_n86, gm_n2788, gm_n2182);
	nor (gm_n2790, gm_n55, in_30, in_29, gm_n2789, gm_n1050);
	nand (gm_n2791, gm_n110, in_12, in_8, gm_n257, gm_n189);
	nor (gm_n2792, gm_n374, in_20, in_16, gm_n2791, gm_n476);
	nand (gm_n2793, gm_n339, gm_n83, in_24, gm_n2792, gm_n263);
	nor (gm_n2794, gm_n2793, gm_n234);
	nand (gm_n2795, gm_n730, gm_n128, gm_n218);
	nor (gm_n2796, gm_n613, in_15, in_11, gm_n2795, gm_n623);
	nand (gm_n2797, gm_n173, gm_n158, gm_n58, gm_n2796, gm_n391);
	nor (gm_n2798, gm_n423, in_31, gm_n54, gm_n2797);
	nor (gm_n2799, gm_n670, in_15, gm_n61, gm_n1723, gm_n398);
	nand (gm_n2800, gm_n513, in_23, gm_n58, gm_n2799, gm_n1042);
	nor (gm_n2801, gm_n618, gm_n55, gm_n54, gm_n2800, gm_n583);
	nor (gm_n2802, gm_n2794, gm_n2790, gm_n2787, gm_n2801, gm_n2798);
	nand (gm_n2803, gm_n731, gm_n71);
	nor (gm_n2804, gm_n188, in_12, in_8, gm_n2803, gm_n237);
	nand (gm_n2805, gm_n103, in_20, gm_n73, gm_n2804, gm_n521);
	nor (gm_n2806, gm_n195, in_28, in_24, gm_n2805, gm_n216);
	nor (gm_n2807, gm_n553, in_16, gm_n63, gm_n1117, gm_n599);
	nand (gm_n2808, gm_n90, gm_n82, in_20, gm_n2807, gm_n263);
	nor (gm_n2809, gm_n214, gm_n85, gm_n83, gm_n2808);
	nor (gm_n2810, gm_n725, in_15, gm_n61, gm_n503, gm_n669);
	nand (gm_n2811, gm_n302, in_23, gm_n58, gm_n2810, gm_n358);
	nor (gm_n2812, gm_n422, gm_n55, gm_n54, gm_n2811, gm_n612);
	nor (gm_n2813, gm_n2812, gm_n2809, gm_n2806);
	nor (gm_n2814, gm_n725, in_15, gm_n61, gm_n822, gm_n363);
	nand (gm_n2815, gm_n296, in_23, gm_n58, gm_n2814, gm_n359);
	nor (gm_n2816, gm_n612, in_31, in_27, gm_n2815, gm_n458);
	nor (gm_n2817, gm_n669, in_15, gm_n61, gm_n1479, gm_n670);
	nand (gm_n2818, gm_n174, gm_n158, in_19, gm_n2817, gm_n334);
	nor (gm_n2819, gm_n423, gm_n55, gm_n54, gm_n2818, gm_n583);
	nand (gm_n2820, gm_n311, gm_n189);
	nor (gm_n2821, gm_n619, gm_n62, in_11, gm_n2820, gm_n425);
	nand (gm_n2822, gm_n77, in_23, gm_n58, gm_n2821, gm_n121);
	nor (gm_n2823, gm_n437, gm_n55, gm_n54, gm_n2822, gm_n458);
	nor (gm_n2824, gm_n2823, gm_n2819, gm_n2816);
	nand (gm_n2825, gm_n2802, gm_n2784, gm_n2781, gm_n2824, gm_n2813);
	nand (gm_n2826, gm_n455, gm_n62, in_11, gm_n2577, gm_n1226);
	nor (gm_n2827, gm_n514, gm_n158, in_19, gm_n2826, gm_n977);
	nand (gm_n2828, gm_n308, in_31, gm_n54, gm_n2827);
	nor (gm_n2829, gm_n93, in_12, gm_n124, gm_n288, gm_n168);
	nand (gm_n2830, gm_n200, in_20, in_16, gm_n2829, gm_n141);
	nor (gm_n2831, gm_n224, gm_n83, in_24, gm_n2830, gm_n411);
	nand (gm_n2832, gm_n2831, gm_n101);
	and (gm_n2833, gm_n123, gm_n62, in_8, gm_n1899, gm_n256);
	nand (gm_n2834, gm_n174, gm_n158, in_19, gm_n2833, gm_n316);
	or (gm_n2835, gm_n57, gm_n55, in_27, gm_n2834, gm_n977);
	nand (gm_n2836, gm_n2835, gm_n2832, gm_n2828);
	nand (gm_n2837, gm_n424, in_15, gm_n61, gm_n792, gm_n426);
	nor (gm_n2838, gm_n131, gm_n158, in_19, gm_n2837, gm_n393);
	nand (gm_n2839, gm_n56, in_31, gm_n54, gm_n2838, gm_n182);
	nand (gm_n2840, gm_n200, in_16, in_12, gm_n887, gm_n110);
	nor (gm_n2841, gm_n197, gm_n82, gm_n76, gm_n2840, gm_n801);
	nand (gm_n2842, gm_n466, gm_n225, in_28, gm_n2841);
	nor (gm_n2843, gm_n669, gm_n93, in_11, gm_n469, gm_n619);
	nand (gm_n2844, gm_n121, in_19, gm_n62, gm_n2843, gm_n130);
	nor (gm_n2845, gm_n183, in_27, gm_n158, gm_n2844, gm_n423);
	nand (gm_n2846, gm_n2845, gm_n55);
	nand (gm_n2847, gm_n2846, gm_n2842, gm_n2839);
	nor (gm_n2848, gm_n2825, gm_n2778, gm_n2775, gm_n2847, gm_n2836);
	nor (gm_n2849, gm_n322, gm_n62, gm_n61, gm_n986, gm_n398);
	nand (gm_n2850, gm_n513, gm_n158, in_19, gm_n2849, gm_n1042);
	nor (gm_n2851, gm_n183, gm_n55, in_27, gm_n2850, gm_n618);
	nor (gm_n2852, gm_n109, gm_n73, gm_n63, gm_n1023, gm_n599);
	nand (gm_n2853, gm_n255, gm_n82, gm_n76, gm_n2852, gm_n477);
	nor (gm_n2854, gm_n224, gm_n185, gm_n83, gm_n2853);
	nor (gm_n2855, gm_n282, in_15, gm_n124, gm_n991, gm_n384);
	nand (gm_n2856, gm_n77, gm_n158, gm_n58, gm_n2855, gm_n121);
	nor (gm_n2857, gm_n423, gm_n55, in_27, gm_n2856, gm_n458);
	nor (gm_n2858, gm_n2857, gm_n2854, gm_n2851);
	nor (gm_n2859, gm_n197, gm_n76, in_16, gm_n2791, gm_n188);
	nand (gm_n2860, gm_n84, gm_n83, in_24, gm_n2859, gm_n192);
	nor (gm_n2861, gm_n2860, gm_n195);
	nor (gm_n2862, gm_n398, gm_n62, in_11, gm_n2682, gm_n619);
	nand (gm_n2863, gm_n121, gm_n158, gm_n58, gm_n2862, gm_n513);
	nor (gm_n2864, gm_n57, gm_n55, in_27, gm_n2863, gm_n512);
	nor (gm_n2865, gm_n92, gm_n73, in_12, gm_n2032, gm_n374);
	nand (gm_n2866, gm_n103, in_24, in_20, gm_n2865, gm_n477);
	nor (gm_n2867, gm_n774, gm_n185, gm_n83, gm_n2866);
	nor (gm_n2868, gm_n2867, gm_n2864, gm_n2861);
	nand (gm_n2869, gm_n2848, gm_n2772, gm_n2769, gm_n2868, gm_n2858);
	or (gm_n2870, gm_n168, gm_n152, in_8);
	nor (gm_n2871, gm_n374, in_16, in_12, gm_n2870, gm_n282);
	and (gm_n2872, gm_n164, in_24, gm_n76, gm_n2871, gm_n227);
	nand (gm_n2873, gm_n137, gm_n102, in_28, gm_n2872);
	nand (gm_n2874, gm_n176, gm_n73, gm_n63, gm_n2096, gm_n340);
	nor (gm_n2875, gm_n411, gm_n82, in_20, gm_n2874, gm_n412);
	nand (gm_n2876, gm_n466, gm_n81, in_28, gm_n2875);
	or (gm_n2877, gm_n109, in_16, in_12, gm_n1519, gm_n288);
	nor (gm_n2878, gm_n197, in_24, in_20, gm_n2877, gm_n411);
	nand (gm_n2879, gm_n225, gm_n102, gm_n83, gm_n2878);
	nand (gm_n2880, gm_n2879, gm_n2876, gm_n2873);
	and (gm_n2881, gm_n66, gm_n198, in_8, gm_n208, gm_n218);
	nor (gm_n2882, in_13, gm_n63, in_11);
	nand (gm_n2883, gm_n486, in_18, in_14, gm_n2882, gm_n2881);
	nor (gm_n2884, gm_n638, in_26, gm_n87, gm_n2883, gm_n1895);
	nand (gm_n2885, gm_n492, gm_n55, gm_n100, gm_n2884);
	or (gm_n2886, gm_n188, in_16, in_12, gm_n1719, gm_n237);
	nor (gm_n2887, gm_n108, gm_n82, in_20, gm_n2886, gm_n801);
	nand (gm_n2888, gm_n225, gm_n186, gm_n83, gm_n2887);
	nand (gm_n2889, gm_n126, gm_n62, in_11, gm_n1676, gm_n313);
	nor (gm_n2890, gm_n303, in_23, in_19, gm_n2889, gm_n431);
	nand (gm_n2891, gm_n60, gm_n55, in_27, gm_n2890, gm_n511);
	nand (gm_n2892, gm_n2891, gm_n2888, gm_n2885);
	nor (gm_n2893, gm_n2869, gm_n2765, gm_n2762, gm_n2892, gm_n2880);
	and (gm_n2894, gm_n167, in_16, gm_n63, gm_n1491, gm_n176);
	nand (gm_n2895, gm_n90, gm_n82, in_20, gm_n2894, gm_n227);
	nor (gm_n2896, gm_n216, gm_n214, in_28, gm_n2895);
	and (gm_n2897, gm_n797, gm_n62, gm_n61, gm_n1226, gm_n544);
	nand (gm_n2898, gm_n174, gm_n158, gm_n58, gm_n2897, gm_n334);
	nor (gm_n2899, gm_n422, in_31, gm_n54, gm_n2898, gm_n675);
	and (gm_n2900, gm_n142, gm_n63, in_8, gm_n1946, gm_n340);
	nand (gm_n2901, gm_n90, gm_n76, gm_n73, gm_n2900, gm_n103);
	nor (gm_n2902, gm_n248, gm_n83, gm_n82, gm_n2901, gm_n195);
	nor (gm_n2903, gm_n2902, gm_n2899, gm_n2896);
	nor (gm_n2904, gm_n432, gm_n58, in_15, gm_n2256, gm_n331);
	nand (gm_n2905, gm_n182, gm_n54, in_23, gm_n2904, gm_n358);
	nor (gm_n2906, gm_n2905, gm_n357, gm_n55);
	nor (gm_n2907, gm_n154, in_16, in_12, gm_n1046, gm_n374);
	nand (gm_n2908, gm_n192, in_24, gm_n76, gm_n2907, gm_n477);
	nor (gm_n2909, gm_n224, gm_n234, gm_n83, gm_n2908);
	and (gm_n2910, gm_n698, in_15, gm_n61, gm_n544, gm_n394);
	nand (gm_n2911, gm_n334, gm_n158, gm_n58, gm_n2910, gm_n455);
	nor (gm_n2912, gm_n357, gm_n55, in_27, gm_n2911, gm_n977);
	nor (gm_n2913, gm_n2912, gm_n2909, gm_n2906);
	nand (gm_n2914, gm_n2893, gm_n2759, gm_n2756, gm_n2913, gm_n2903);
	nor (gm_n2915, gm_n670, gm_n62, gm_n61, gm_n758, gm_n623);
	nand (gm_n2916, gm_n513, gm_n158, in_19, gm_n2915, gm_n1042);
	nor (gm_n2917, gm_n423, gm_n55, in_27, gm_n2916, gm_n583);
	or (gm_n2918, gm_n154, in_12, gm_n124, gm_n345, gm_n168);
	or (gm_n2919, gm_n143, gm_n76, in_16, gm_n2918, gm_n463);
	or (gm_n2920, gm_n216, gm_n83, gm_n82, gm_n2919, gm_n566);
	nor (gm_n2921, gm_n2920, gm_n195);
	and (gm_n2922, gm_n797, in_15, gm_n61, gm_n699, gm_n622);
	and (gm_n2923, gm_n121, gm_n158, in_19, gm_n2922, gm_n334);
	and (gm_n2924, gm_n56, gm_n55, gm_n54, gm_n2923, gm_n459);
	nor (gm_n2925, gm_n2924, gm_n2921, gm_n2917);
	not (gm_n2926, gm_n2925);
	nor (gm_n2927, gm_n111, in_12, in_8, gm_n1038, gm_n236);
	nand (gm_n2928, gm_n235, in_20, in_16, gm_n2927, gm_n263);
	nor (gm_n2929, gm_n185, in_28, in_24, gm_n2928, gm_n262);
	or (gm_n2930, gm_n2914, gm_n2753, gm_n2750, gm_n2929, gm_n2926);
	not (gm_n2931, t_2);
	nor (gm_n2932, gm_n374, gm_n73, in_12, gm_n1979, gm_n282);
	nand (gm_n2933, gm_n88, gm_n82, gm_n76, gm_n2932, gm_n477);
	nor (gm_n2934, gm_n262, gm_n214, gm_n83, gm_n2933);
	and (gm_n2935, gm_n797, in_15, in_11, gm_n332, gm_n123);
	nand (gm_n2936, gm_n455, in_23, in_19, gm_n2935, gm_n513);
	nor (gm_n2937, gm_n57, in_31, in_27, gm_n2936, gm_n977);
	nor (gm_n2938, gm_n111, gm_n73, in_12, gm_n238, gm_n188);
	and (gm_n2939, gm_n263, in_24, gm_n76, gm_n2938, gm_n477);
	and (gm_n2940, gm_n367, gm_n225, gm_n83, gm_n2939);
	and (gm_n2941, gm_n995, in_15, in_11, gm_n2581, gm_n1226);
	nand (gm_n2942, gm_n130, in_23, in_19, gm_n2941, gm_n174);
	or (gm_n2943, gm_n422, gm_n55, in_27, gm_n2942, gm_n437);
	or (gm_n2944, gm_n179, in_20, gm_n73, gm_n522, gm_n188);
	nor (gm_n2945, gm_n224, gm_n83, gm_n82, gm_n2944, gm_n520);
	nand (gm_n2946, gm_n2945, gm_n213);
	nor (gm_n2947, gm_n374, gm_n73, gm_n63, gm_n2070, gm_n237);
	nand (gm_n2948, gm_n205, in_24, in_20, gm_n2947, gm_n477);
	nor (gm_n2949, gm_n216, gm_n195, gm_n83, gm_n2948);
	nand (gm_n2950, gm_n218, in_12, in_8, gm_n731, gm_n153);
	nor (gm_n2951, gm_n197, in_20, gm_n73, gm_n2950, gm_n374);
	and (gm_n2952, gm_n88, gm_n83, gm_n82, gm_n2951, gm_n367);
	and (gm_n2953, gm_n2952, gm_n81);
	and (gm_n2954, gm_n128, gm_n63, in_8, gm_n310, gm_n242);
	and (gm_n2955, gm_n446, gm_n76, gm_n73, gm_n2954, gm_n235);
	and (gm_n2956, gm_n339, gm_n83, gm_n82, gm_n2955, gm_n263);
	and (gm_n2957, gm_n2956, gm_n101);
	nand (gm_n2958, gm_n167, gm_n63, in_8, gm_n1133, gm_n176);
	or (gm_n2959, gm_n104, in_20, gm_n73, gm_n2958, gm_n108);
	nor (gm_n2960, gm_n248, gm_n83, gm_n82, gm_n2959, gm_n214);
	and (gm_n2961, gm_n71, in_12, in_8, gm_n594, gm_n167);
	and (gm_n2962, gm_n90, gm_n76, gm_n73, gm_n2961, gm_n200);
	and (gm_n2963, gm_n102, gm_n83, gm_n82, gm_n2962, gm_n217);
	and (gm_n2964, gm_n2963, gm_n81);
	nand (gm_n2965, gm_n153, gm_n73, gm_n63, gm_n1499, gm_n166);
	or (gm_n2966, gm_n801, in_24, in_20, gm_n2965, gm_n476);
	nor (gm_n2967, gm_n216, gm_n234, in_28, gm_n2966);
	or (gm_n2968, gm_n433, in_15, in_11, gm_n991, gm_n874);
	nor (gm_n2969, gm_n335, in_23, in_19, gm_n2968, gm_n456);
	and (gm_n2970, gm_n305, gm_n55, gm_n54, gm_n2969, gm_n511);
	nor (gm_n2971, gm_n282, in_15, gm_n124, gm_n384, gm_n363);
	nand (gm_n2972, gm_n77, in_23, gm_n58, gm_n2971, gm_n359);
	nor (gm_n2973, gm_n583, gm_n55, in_27, gm_n2972, gm_n838);
	nor (gm_n2974, gm_n249, gm_n73, gm_n63, gm_n2070, gm_n92);
	nand (gm_n2975, gm_n107, gm_n82, gm_n76, gm_n2974, gm_n192);
	nor (gm_n2976, gm_n684, gm_n140, in_28, gm_n2975);
	and (gm_n2977, gm_n200, in_12, gm_n124, gm_n1899, gm_n242);
	nand (gm_n2978, gm_n141, in_20, in_16, gm_n2977, gm_n192);
	nor (gm_n2979, gm_n214, in_28, gm_n82, gm_n2978, gm_n774);
	nand (gm_n2980, gm_n200, in_16, gm_n63, gm_n201, gm_n153);
	or (gm_n2981, gm_n187, in_24, in_20, gm_n2980, gm_n566);
	nor (gm_n2982, gm_n185, gm_n85, gm_n83, gm_n2981);
	or (gm_n2983, gm_n2976, gm_n2973, gm_n2970, gm_n2982, gm_n2979);
	nand (gm_n2984, gm_n110, gm_n73, in_12, gm_n572, gm_n142);
	or (gm_n2985, gm_n89, gm_n82, in_20, gm_n2984, gm_n412);
	nor (gm_n2986, gm_n214, gm_n248, gm_n83, gm_n2985);
	and (gm_n2987, gm_n207, in_16, in_12, gm_n1706, gm_n228);
	nand (gm_n2988, gm_n217, in_24, in_20, gm_n2987, gm_n477);
	nor (gm_n2989, gm_n684, gm_n368, gm_n83, gm_n2988);
	or (gm_n2990, gm_n669, gm_n62, gm_n61, gm_n1209, gm_n619);
	nor (gm_n2991, gm_n331, gm_n158, in_19, gm_n2990, gm_n335);
	and (gm_n2992, gm_n305, gm_n55, gm_n54, gm_n2991, gm_n674);
	or (gm_n2993, gm_n2992, gm_n2989, gm_n2986);
	or (gm_n2994, gm_n154, gm_n73, in_12, gm_n776, gm_n188);
	or (gm_n2995, gm_n108, in_24, gm_n76, gm_n2994, gm_n801);
	nor (gm_n2996, gm_n684, gm_n224, gm_n83, gm_n2995);
	or (gm_n2997, gm_n125, gm_n62, gm_n61, gm_n2491, gm_n623);
	or (gm_n2998, gm_n331, gm_n158, in_19, gm_n2997, gm_n317);
	nor (gm_n2999, gm_n618, in_31, gm_n54, gm_n2998, gm_n977);
	or (gm_n3000, gm_n122, gm_n158, in_19, gm_n1615, gm_n335);
	nor (gm_n3001, gm_n583, gm_n55, in_27, gm_n3000, gm_n838);
	or (gm_n3002, gm_n3001, gm_n2999, gm_n2996);
	or (gm_n3003, gm_n2983, gm_n2967, gm_n2964, gm_n3002, gm_n2993);
	or (gm_n3004, gm_n669, in_15, in_11, gm_n1272, gm_n322);
	or (gm_n3005, gm_n796, in_23, gm_n58, gm_n3004, gm_n317);
	nor (gm_n3006, gm_n512, gm_n55, gm_n54, gm_n3005, gm_n618);
	nand (gm_n3007, gm_n142, gm_n73, gm_n63, gm_n2555, gm_n228);
	or (gm_n3008, gm_n187, gm_n82, gm_n76, gm_n3007, gm_n411);
	nor (gm_n3009, gm_n684, gm_n774, in_28, gm_n3008);
	nand (gm_n3010, gm_n65, gm_n58, gm_n62, gm_n1990, gm_n174);
	or (gm_n3011, gm_n335, gm_n54, gm_n158, gm_n3010, gm_n977);
	nor (gm_n3012, gm_n3011, gm_n618, gm_n55);
	or (gm_n3013, gm_n3012, gm_n3009, gm_n3006);
	nor (gm_n3014, gm_n432, in_15, in_11, gm_n2589, gm_n433);
	nand (gm_n3015, gm_n173, in_23, in_19, gm_n3014, gm_n455);
	nor (gm_n3016, gm_n512, gm_n55, gm_n54, gm_n3015, gm_n437);
	or (gm_n3017, gm_n154, gm_n73, gm_n63, gm_n2245, gm_n374);
	or (gm_n3018, gm_n108, in_24, in_20, gm_n3017, gm_n520);
	nor (gm_n3019, gm_n214, gm_n224, gm_n83, gm_n3018);
	or (gm_n3020, gm_n395, in_15, gm_n61, gm_n554, gm_n425);
	or (gm_n3021, gm_n303, in_23, in_19, gm_n3020, gm_n335);
	nor (gm_n3022, gm_n618, in_31, gm_n54, gm_n3021, gm_n458);
	or (gm_n3023, gm_n3022, gm_n3019, gm_n3016);
	or (gm_n3024, gm_n3003, gm_n2960, gm_n2957, gm_n3023, gm_n3013);
	nor (gm_n3025, gm_n447, in_12, in_8, gm_n178, gm_n154);
	and (gm_n3026, gm_n166, gm_n76, gm_n73, gm_n3025, gm_n477);
	and (gm_n3027, gm_n186, in_28, gm_n82, gm_n3026, gm_n255);
	and (gm_n3028, gm_n3027, gm_n496);
	nor (gm_n3029, gm_n152, gm_n63, gm_n124, gm_n288, gm_n271);
	and (gm_n3030, gm_n142, in_20, gm_n73, gm_n3029, gm_n164);
	and (gm_n3031, gm_n139, gm_n83, in_24, gm_n3030, gm_n205);
	and (gm_n3032, gm_n3031, gm_n629);
	nor (gm_n3033, gm_n249, in_16, gm_n63, gm_n2870, gm_n237);
	nand (gm_n3034, gm_n107, gm_n82, in_20, gm_n3033, gm_n263);
	nor (gm_n3035, gm_n214, gm_n85, in_28, gm_n3034);
	or (gm_n3036, gm_n3035, gm_n3032, gm_n3028);
	nand (gm_n3037, gm_n199, gm_n73, gm_n63, gm_n1590, gm_n207);
	or (gm_n3038, gm_n801, gm_n82, in_20, gm_n3037, gm_n476);
	nor (gm_n3039, gm_n195, gm_n224, in_28, gm_n3038);
	nand (gm_n3040, gm_n995, gm_n62, gm_n61, gm_n2142, gm_n698);
	or (gm_n3041, gm_n335, in_23, in_19, gm_n3040, gm_n360);
	nor (gm_n3042, gm_n57, gm_n55, in_27, gm_n3041, gm_n512);
	nand (gm_n3043, gm_n150, in_16, gm_n63, gm_n1740, gm_n256);
	or (gm_n3044, gm_n187, gm_n82, in_20, gm_n3043, gm_n520);
	nor (gm_n3045, gm_n226, gm_n224, gm_n83, gm_n3044);
	or (gm_n3046, gm_n3045, gm_n3042, gm_n3039);
	nor (gm_n3047, gm_n3024, gm_n2953, gm_n2949, gm_n3046, gm_n3036);
	and (gm_n3048, gm_n71, gm_n63, in_8, gm_n208, gm_n167);
	and (gm_n3049, gm_n150, gm_n76, gm_n73, gm_n3048, gm_n477);
	and (gm_n3050, gm_n102, in_28, in_24, gm_n3049, gm_n263);
	and (gm_n3051, gm_n3050, gm_n101);
	nor (gm_n3052, gm_n249, in_16, gm_n63, gm_n558, gm_n154);
	nand (gm_n3053, gm_n88, in_24, in_20, gm_n3052, gm_n235);
	nor (gm_n3054, gm_n479, gm_n774, in_28, gm_n3053);
	nor (gm_n3055, gm_n664, gm_n62, in_11, gm_n991, gm_n874);
	and (gm_n3056, gm_n296, gm_n158, gm_n58, gm_n3055, gm_n455);
	and (gm_n3057, gm_n305, in_31, in_27, gm_n3056, gm_n511);
	nor (gm_n3058, gm_n3057, gm_n3054, gm_n3051);
	and (gm_n3059, gm_n189, gm_n63, in_8, gm_n257, gm_n256);
	and (gm_n3060, gm_n446, in_20, gm_n73, gm_n3059, gm_n270);
	and (gm_n3061, gm_n217, gm_n83, gm_n82, gm_n3060, gm_n339);
	and (gm_n3062, gm_n3061, gm_n496);
	nor (gm_n3063, in_21, gm_n76, in_19);
	and (gm_n3064, gm_n1893, in_22, gm_n106, gm_n3063, gm_n2464);
	nand (gm_n3065, gm_n3064, gm_n639, in_26);
	nor (gm_n3066, gm_n2446, gm_n55, in_30, gm_n3065);
	nor (gm_n3067, gm_n725, in_15, gm_n61, gm_n1805, gm_n669);
	nand (gm_n3068, gm_n121, in_23, gm_n58, gm_n3067, gm_n358);
	nor (gm_n3069, gm_n1200, in_31, in_27, gm_n3068, gm_n612);
	nor (gm_n3070, gm_n3069, gm_n3066, gm_n3062);
	nand (gm_n3071, gm_n3047, gm_n2946, gm_n2943, gm_n3070, gm_n3058);
	nand (gm_n3072, gm_n207, gm_n73, in_12, gm_n549, gm_n256);
	nor (gm_n3073, gm_n89, gm_n82, gm_n76, gm_n3072, gm_n476);
	nand (gm_n3074, gm_n225, gm_n139, gm_n83, gm_n3073);
	nand (gm_n3075, gm_n446, gm_n73, in_12, gm_n1740, gm_n242);
	nor (gm_n3076, gm_n630, gm_n82, gm_n76, gm_n3075, gm_n412);
	nand (gm_n3077, gm_n496, gm_n102, in_28, gm_n3076);
	nand (gm_n3078, gm_n167, gm_n73, in_12, gm_n230, gm_n207);
	nor (gm_n3079, gm_n206, in_24, in_20, gm_n3078, gm_n522);
	nand (gm_n3080, gm_n137, gm_n102, gm_n83, gm_n3079);
	nand (gm_n3081, gm_n3080, gm_n3077, gm_n3074);
	nand (gm_n3082, gm_n153, in_16, in_12, gm_n1574, gm_n207);
	nor (gm_n3083, gm_n463, in_24, gm_n76, gm_n3082, gm_n630);
	nand (gm_n3084, gm_n466, gm_n196, gm_n83, gm_n3083);
	or (gm_n3085, gm_n92, gm_n73, gm_n63, gm_n2046, gm_n143);
	nor (gm_n3086, gm_n165, in_24, in_20, gm_n3085, gm_n801);
	nand (gm_n3087, gm_n215, gm_n213, in_28, gm_n3086);
	nand (gm_n3088, gm_n1630, gm_n65, gm_n62);
	nor (gm_n3089, gm_n331, gm_n158, in_19, gm_n3088, gm_n317);
	nand (gm_n3090, gm_n60, gm_n55, gm_n54, gm_n3089, gm_n674);
	nand (gm_n3091, gm_n3090, gm_n3087, gm_n3084);
	or (gm_n3092, gm_n3071, gm_n2940, gm_n2937, gm_n3091, gm_n3081);
	and (gm_n3093, gm_n199, gm_n65, in_15, gm_n1706, gm_n455);
	nand (gm_n3094, gm_n60, in_23, gm_n58, gm_n3093, gm_n173);
	nor (gm_n3095, gm_n423, in_31, in_27, gm_n3094);
	nor (gm_n3096, gm_n249, gm_n63, gm_n124, gm_n1164, gm_n282);
	and (gm_n3097, gm_n235, gm_n76, in_16, gm_n3096, gm_n263);
	and (gm_n3098, gm_n81, in_28, in_24, gm_n3097, gm_n84);
	and (gm_n3099, gm_n142, in_16, in_12, gm_n572, gm_n228);
	and (gm_n3100, gm_n227, in_24, in_20, gm_n3099, gm_n235);
	and (gm_n3101, gm_n367, gm_n101, gm_n83, gm_n3100);
	nor (gm_n3102, gm_n3101, gm_n3098, gm_n3095);
	not (gm_n3103, gm_n3102);
	nand (gm_n3104, gm_n731, gm_n144, gm_n124);
	nor (gm_n3105, gm_n111, gm_n73, in_12, gm_n3104, gm_n177);
	and (gm_n3106, gm_n192, in_24, in_20, gm_n3105, gm_n235);
	and (gm_n3107, gm_n196, gm_n84, gm_n83, gm_n3106);
	or (gm_n3108, gm_n3092, gm_n2934, gm_n2931, gm_n3107, gm_n3103);
	nand (gm_n3109, gm_n3108, gm_n2930);
	not (gm_n3110, t_1);
	or (gm_n3111, gm_n303, in_19, in_15, gm_n623, gm_n579);
	or (gm_n3112, gm_n422, in_27, in_23, gm_n3111, gm_n431);
	nor (gm_n3113, gm_n3112, gm_n838, gm_n55);
	nand (gm_n3114, gm_n66, in_9, gm_n124, gm_n703, gm_n127);
	or (gm_n3115, gm_n122, gm_n62, gm_n61, gm_n3114, gm_n314);
	or (gm_n3116, gm_n452, gm_n158, gm_n58, gm_n3115, gm_n458);
	nor (gm_n3117, gm_n423, in_31, gm_n54, gm_n3116);
	nor (gm_n3118, gm_n109, gm_n73, in_12, gm_n2327, gm_n237);
	and (gm_n3119, gm_n141, gm_n82, in_20, gm_n3118, gm_n217);
	and (gm_n3120, gm_n137, gm_n84, gm_n83, gm_n3119);
	nand (gm_n3121, gm_n426, in_15, in_11, gm_n699, gm_n730);
	nor (gm_n3122, gm_n331, gm_n158, in_19, gm_n3121, gm_n317);
	nand (gm_n3123, gm_n305, gm_n55, in_27, gm_n3122, gm_n337);
	not (gm_n3124, gm_n1679);
	nand (gm_n3125, gm_n76, in_19, gm_n106);
	or (gm_n3126, gm_n534, gm_n86, in_17, gm_n3125, gm_n1677);
	nor (gm_n3127, gm_n160, gm_n80, in_25, gm_n3126, gm_n3124);
	nand (gm_n3128, gm_n3127, in_31, in_30);
	nand (gm_n3129, gm_n199, gm_n73, gm_n63, gm_n220, gm_n207);
	or (gm_n3130, gm_n801, gm_n82, in_20, gm_n3129, gm_n412);
	nor (gm_n3131, gm_n774, gm_n195, in_28, gm_n3130);
	nand (gm_n3132, gm_n142, gm_n73, gm_n63, gm_n900, gm_n153);
	or (gm_n3133, gm_n206, gm_n82, in_20, gm_n3132, gm_n476);
	nor (gm_n3134, gm_n368, gm_n226, gm_n83, gm_n3133);
	nand (gm_n3135, gm_n123, gm_n62, gm_n61, gm_n1400, gm_n300);
	nor (gm_n3136, gm_n317, in_23, in_19, gm_n3135, gm_n613);
	nand (gm_n3137, gm_n134, in_31, gm_n54, gm_n3136, gm_n511);
	and (gm_n3138, gm_n176, gm_n73, gm_n63, gm_n2514, gm_n340);
	nand (gm_n3139, gm_n227, in_24, in_20, gm_n3138, gm_n270);
	or (gm_n3140, gm_n195, gm_n248, gm_n83, gm_n3139);
	nor (gm_n3141, gm_n111, gm_n73, in_12, gm_n1100, gm_n177);
	nand (gm_n3142, gm_n205, in_24, gm_n76, gm_n3141, gm_n235);
	nor (gm_n3143, gm_n368, gm_n185, in_28, gm_n3142);
	and (gm_n3144, gm_n200, gm_n73, in_12, gm_n2567, gm_n110);
	nand (gm_n3145, gm_n90, in_24, in_20, gm_n3144, gm_n103);
	nor (gm_n3146, gm_n684, gm_n774, gm_n83, gm_n3145);
	nand (gm_n3147, gm_n150, gm_n73, gm_n63, gm_n900, gm_n340);
	nor (gm_n3148, gm_n104, in_24, in_20, gm_n3147, gm_n522);
	nand (gm_n3149, gm_n496, gm_n139, gm_n83, gm_n3148);
	and (gm_n3150, gm_n455, gm_n340, gm_n62, gm_n1706, gm_n622);
	nand (gm_n3151, gm_n173, gm_n158, gm_n58, gm_n3150, gm_n182);
	or (gm_n3152, gm_n618, gm_n55, in_27, gm_n3151);
	nor (gm_n3153, gm_n322, gm_n62, gm_n61, gm_n434, gm_n398);
	and (gm_n3154, gm_n77, gm_n158, gm_n58, gm_n3153, gm_n455);
	nand (gm_n3155, gm_n134, in_31, in_27, gm_n3154, gm_n674);
	or (gm_n3156, gm_n109, gm_n73, gm_n63, gm_n952, gm_n282);
	nor (gm_n3157, gm_n520, in_24, in_20, gm_n3156, gm_n522);
	nand (gm_n3158, gm_n225, gm_n215, in_28, gm_n3157);
	nor (gm_n3159, gm_n188, gm_n73, gm_n63, gm_n288, gm_n250);
	and (gm_n3160, gm_n217, gm_n82, in_20, gm_n3159, gm_n270);
	nand (gm_n3161, gm_n102, gm_n81, in_28, gm_n3160);
	nand (gm_n3162, gm_n3155, gm_n3152, gm_n3149, gm_n3161, gm_n3158);
	and (gm_n3163, gm_n300, in_15, gm_n61, gm_n1791, gm_n931);
	nand (gm_n3164, gm_n121, gm_n158, gm_n58, gm_n3163, gm_n130);
	or (gm_n3165, gm_n57, in_31, in_27, gm_n3164, gm_n977);
	nand (gm_n3166, gm_n123, gm_n62, in_11, gm_n2128, gm_n359);
	nor (gm_n3167, gm_n431, in_23, gm_n58, gm_n3166, gm_n977);
	nand (gm_n3168, gm_n337, in_31, in_27, gm_n3167);
	and (gm_n3169, gm_n394, gm_n127, in_11, gm_n622, gm_n588);
	nand (gm_n3170, gm_n130, in_19, in_15, gm_n3169, gm_n302);
	nor (gm_n3171, gm_n57, in_27, gm_n158, gm_n3170, gm_n422);
	nand (gm_n3172, gm_n3171, in_31);
	nand (gm_n3173, gm_n3172, gm_n3168, gm_n3165);
	nand (gm_n3174, gm_n703, gm_n127, in_8);
	or (gm_n3175, gm_n599, gm_n73, gm_n63, gm_n3174, gm_n188);
	nor (gm_n3176, gm_n801, in_24, in_20, gm_n3175, gm_n476);
	nand (gm_n3177, gm_n102, gm_n101, in_28, gm_n3176);
	and (gm_n3178, gm_n110, in_16, in_12, gm_n567, gm_n142);
	and (gm_n3179, gm_n205, gm_n82, gm_n76, gm_n3178, gm_n477);
	nand (gm_n3180, gm_n215, gm_n81, in_28, gm_n3179);
	nand (gm_n3181, gm_n199, gm_n73, gm_n63, gm_n2486, gm_n166);
	nor (gm_n3182, gm_n566, gm_n82, in_20, gm_n3181, gm_n476);
	nand (gm_n3183, gm_n367, gm_n101, in_28, gm_n3182);
	nand (gm_n3184, gm_n3183, gm_n3180, gm_n3177);
	nor (gm_n3185, gm_n3162, gm_n3146, gm_n3143, gm_n3184, gm_n3173);
	nor (gm_n3186, gm_n432, gm_n62, in_11, gm_n1252, gm_n125);
	nand (gm_n3187, gm_n77, in_23, gm_n58, gm_n3186, gm_n1042);
	nor (gm_n3188, gm_n183, in_31, in_27, gm_n3187, gm_n618);
	nor (gm_n3189, gm_n109, in_16, in_12, gm_n631, gm_n599);
	nand (gm_n3190, gm_n164, in_24, in_20, gm_n3189, gm_n192);
	nor (gm_n3191, gm_n248, gm_n138, gm_n83, gm_n3190);
	nor (gm_n3192, gm_n236, gm_n73, gm_n63, gm_n1296, gm_n237);
	nand (gm_n3193, gm_n103, in_24, gm_n76, gm_n3192, gm_n270);
	nor (gm_n3194, gm_n774, gm_n226, in_28, gm_n3193);
	nor (gm_n3195, gm_n3194, gm_n3191, gm_n3188);
	nor (gm_n3196, gm_n236, in_20, in_16, gm_n1088, gm_n522);
	nand (gm_n3197, gm_n205, gm_n83, in_24, gm_n3196, gm_n215);
	nor (gm_n3198, gm_n3197, gm_n195);
	nor (gm_n3199, gm_n111, gm_n73, in_12, gm_n1168, gm_n553);
	nand (gm_n3200, gm_n88, in_24, in_20, gm_n3199, gm_n107);
	nor (gm_n3201, gm_n684, gm_n85, gm_n83, gm_n3200);
	or (gm_n3202, gm_n599, gm_n63, in_8, gm_n345, gm_n277);
	nor (gm_n3203, gm_n187, gm_n76, gm_n73, gm_n3202, gm_n553);
	nand (gm_n3204, gm_n263, gm_n83, in_24, gm_n3203, gm_n367);
	nor (gm_n3205, gm_n3204, gm_n185);
	nor (gm_n3206, gm_n3205, gm_n3201, gm_n3198);
	nand (gm_n3207, gm_n3185, gm_n3140, gm_n3137, gm_n3206, gm_n3195);
	nand (gm_n3208, gm_n65, in_15, gm_n61, gm_n1938, gm_n797);
	or (gm_n3209, gm_n297, gm_n158, gm_n58, gm_n3208, gm_n360);
	nor (gm_n3210, gm_n1200, gm_n55, in_27, gm_n3209, gm_n618);
	and (gm_n3211, gm_n394, gm_n264, in_11, gm_n502);
	and (gm_n3212, gm_n302, in_19, in_15, gm_n3211, gm_n698);
	and (gm_n3213, gm_n391, in_27, in_23, gm_n3212, gm_n513);
	and (gm_n3214, gm_n3213, gm_n438, in_31);
	nand (gm_n3215, gm_n142, in_16, gm_n63, gm_n1904, gm_n153);
	or (gm_n3216, gm_n520, in_24, in_20, gm_n3215, gm_n463);
	nor (gm_n3217, gm_n684, gm_n224, in_28, gm_n3216);
	or (gm_n3218, gm_n3217, gm_n3214, gm_n3210);
	nand (gm_n3219, gm_n150, in_16, in_12, gm_n866, gm_n167);
	or (gm_n3220, gm_n411, gm_n82, in_20, gm_n3219, gm_n522);
	nor (gm_n3221, gm_n85, gm_n234, gm_n83, gm_n3220);
	or (gm_n3222, gm_n116, gm_n63, in_8, gm_n288, gm_n229);
	nor (gm_n3223, gm_n109, in_20, gm_n73, gm_n3222, gm_n463);
	nand (gm_n3224, gm_n103, in_28, gm_n82, gm_n3223, gm_n139);
	nor (gm_n3225, gm_n3224, gm_n185);
	nand (gm_n3226, gm_n207, gm_n76, gm_n73, gm_n2829, gm_n270);
	or (gm_n3227, gm_n566, gm_n83, gm_n82, gm_n3226, gm_n368);
	nor (gm_n3228, gm_n3227, gm_n195);
	or (gm_n3229, gm_n3228, gm_n3225, gm_n3221);
	nor (gm_n3230, gm_n3207, gm_n3134, gm_n3131, gm_n3229, gm_n3218);
	or (gm_n3231, gm_n249, gm_n73, gm_n63, gm_n2032, gm_n237);
	or (gm_n3232, gm_n801, gm_n82, in_20, gm_n3231, gm_n412);
	nor (gm_n3233, gm_n85, gm_n234, in_28, gm_n3232);
	or (gm_n3234, gm_n303, in_23, gm_n58, gm_n3088, gm_n335);
	nor (gm_n3235, gm_n422, in_31, in_27, gm_n3234, gm_n423);
	or (gm_n3236, gm_n188, gm_n73, gm_n63, gm_n3174, gm_n352);
	or (gm_n3237, gm_n104, gm_n82, in_20, gm_n3236, gm_n463);
	nor (gm_n3238, gm_n774, gm_n214, in_28, gm_n3237);
	nor (gm_n3239, gm_n3238, gm_n3235, gm_n3233);
	or (gm_n3240, gm_n374, gm_n63, gm_n124, gm_n2820, gm_n352);
	or (gm_n3241, gm_n89, gm_n76, gm_n73, gm_n3240, gm_n165);
	nor (gm_n3242, gm_n138, gm_n83, in_24, gm_n3241, gm_n140);
	nor (gm_n3243, gm_n143, in_16, gm_n63, gm_n1117, gm_n352);
	nand (gm_n3244, gm_n227, in_24, in_20, gm_n3243, gm_n521);
	nor (gm_n3245, gm_n140, gm_n138, gm_n83, gm_n3244);
	nor (gm_n3246, gm_n146, gm_n62, gm_n61, gm_n991, gm_n395);
	and (gm_n3247, gm_n174, in_23, gm_n58, gm_n3246, gm_n358);
	and (gm_n3248, gm_n459, in_31, gm_n54, gm_n3247, gm_n674);
	nor (gm_n3249, gm_n3248, gm_n3245, gm_n3242);
	nand (gm_n3250, gm_n3230, gm_n3128, gm_n3123, gm_n3249, gm_n3239);
	nor (gm_n3251, gm_n352, gm_n63, in_8, gm_n383, gm_n2141);
	nand (gm_n3252, gm_n446, in_20, in_16, gm_n3251, gm_n521);
	nor (gm_n3253, gm_n85, gm_n83, gm_n82, gm_n3252, gm_n104);
	nand (gm_n3254, gm_n3253, gm_n101);
	nor (gm_n3255, gm_n314, gm_n154, gm_n62, gm_n2070, gm_n613);
	nand (gm_n3256, gm_n60, in_23, in_19, gm_n3255, gm_n130);
	or (gm_n3257, gm_n423, gm_n55, in_27, gm_n3256);
	nor (gm_n3258, gm_n154, in_12, gm_n124, gm_n345, gm_n298);
	nand (gm_n3259, gm_n150, gm_n76, gm_n73, gm_n3258, gm_n521);
	nor (gm_n3260, gm_n89, gm_n83, gm_n82, gm_n3259, gm_n262);
	nand (gm_n3261, gm_n3260, gm_n629);
	nand (gm_n3262, gm_n3261, gm_n3257, gm_n3254);
	nand (gm_n3263, gm_n150, gm_n73, gm_n63, gm_n242, gm_n169);
	nor (gm_n3264, gm_n206, in_24, in_20, gm_n3263, gm_n463);
	nand (gm_n3265, gm_n629, gm_n339, gm_n83, gm_n3264);
	nand (gm_n3266, gm_n121, in_19, gm_n62, gm_n2162, gm_n123);
	nor (gm_n3267, gm_n297, in_27, gm_n158, gm_n3266, gm_n422);
	nand (gm_n3268, gm_n3267, gm_n308, in_31);
	nand (gm_n3269, gm_n142, in_16, in_12, gm_n589, gm_n228);
	nor (gm_n3270, gm_n520, in_24, in_20, gm_n3269, gm_n476);
	nand (gm_n3271, gm_n215, gm_n137, in_28, gm_n3270);
	nand (gm_n3272, gm_n3271, gm_n3268, gm_n3265);
	or (gm_n3273, gm_n3250, gm_n3120, gm_n3117, gm_n3272, gm_n3262);
	nor (gm_n3274, gm_n322, in_15, in_11, gm_n1038, gm_n623);
	and (gm_n3275, gm_n77, gm_n158, in_19, gm_n3274, gm_n174);
	and (gm_n3276, gm_n305, in_31, in_27, gm_n3275, gm_n674);
	nor (gm_n3277, gm_n553, in_12, gm_n124, gm_n2803, gm_n599);
	and (gm_n3278, gm_n88, in_20, in_16, gm_n3277, gm_n164);
	and (gm_n3279, gm_n137, in_28, in_24, gm_n3278, gm_n139);
	and (gm_n3280, gm_n110, gm_n73, gm_n63, gm_n2136, gm_n142);
	and (gm_n3281, gm_n235, in_24, gm_n76, gm_n3280, gm_n263);
	and (gm_n3282, gm_n225, gm_n139, gm_n83, gm_n3281);
	nor (gm_n3283, gm_n3282, gm_n3279, gm_n3276);
	not (gm_n3284, gm_n3283);
	nor (gm_n3285, gm_n395, gm_n62, gm_n61, gm_n2491, gm_n425);
	and (gm_n3286, gm_n77, in_23, gm_n58, gm_n3285, gm_n121);
	and (gm_n3287, gm_n134, gm_n55, gm_n54, gm_n3286, gm_n674);
	or (gm_n3288, gm_n3273, gm_n3113, gm_n3110, gm_n3287, gm_n3284);
	not (gm_n3289, t_0);
	and (gm_n3290, gm_n426, in_19, gm_n62, gm_n1999, gm_n455);
	and (gm_n3291, gm_n77, in_27, in_23, gm_n3290, gm_n182);
	and (gm_n3292, gm_n3291, gm_n674, gm_n55);
	and (gm_n3293, gm_n91, gm_n73, gm_n63, gm_n961, gm_n167);
	and (gm_n3294, gm_n227, gm_n82, gm_n76, gm_n3293, gm_n521);
	and (gm_n3295, gm_n215, gm_n137, in_28, gm_n3294);
	nor (gm_n3296, gm_n432, gm_n62, gm_n61, gm_n874, gm_n433);
	and (gm_n3297, gm_n302, in_23, gm_n58, gm_n3296, gm_n358);
	and (gm_n3298, gm_n459, gm_n55, in_27, gm_n3297, gm_n511);
	nor (gm_n3299, gm_n669, in_15, in_11, gm_n664, gm_n321);
	and (gm_n3300, gm_n358, gm_n158, in_19, gm_n3299, gm_n392);
	and (gm_n3301, gm_n60, gm_n55, in_27, gm_n3300, gm_n308);
	nor (gm_n3302, gm_n143, gm_n63, in_8, gm_n1527, gm_n154);
	and (gm_n3303, gm_n164, gm_n76, gm_n73, gm_n3302, gm_n263);
	nand (gm_n3304, gm_n102, gm_n83, in_24, gm_n3303, gm_n496);
	not (gm_n3305, gm_n3304);
	or (gm_n3306, gm_n670, gm_n62, in_11, gm_n1209, gm_n314);
	or (gm_n3307, gm_n303, in_23, in_19, gm_n3306, gm_n335);
	nor (gm_n3308, gm_n57, in_31, gm_n54, gm_n3307, gm_n458);
	nand (gm_n3309, gm_n126, gm_n62, in_11, gm_n2226, gm_n313);
	or (gm_n3310, gm_n796, gm_n158, gm_n58, gm_n3309, gm_n1225);
	nor (gm_n3311, gm_n1200, gm_n55, in_27, gm_n3310, gm_n838);
	nor (gm_n3312, gm_n432, gm_n62, gm_n61, gm_n986, gm_n619);
	nand (gm_n3313, gm_n296, in_23, gm_n58, gm_n3312, gm_n359);
	nor (gm_n3314, gm_n57, in_31, in_27, gm_n3313, gm_n977);
	or (gm_n3315, gm_n432, gm_n62, gm_n61, gm_n1221, gm_n125);
	or (gm_n3316, gm_n297, in_23, in_19, gm_n3315, gm_n393);
	nor (gm_n3317, gm_n423, gm_n55, in_27, gm_n3316, gm_n977);
	nor (gm_n3318, gm_n432, gm_n62, gm_n61, gm_n1259, gm_n670);
	nand (gm_n3319, gm_n296, in_23, gm_n58, gm_n3318, gm_n1042);
	nor (gm_n3320, gm_n57, in_31, in_27, gm_n3319, gm_n1112);
	or (gm_n3321, gm_n669, in_15, gm_n61, gm_n2381, gm_n360);
	or (gm_n3322, gm_n452, gm_n158, gm_n58, gm_n3321, gm_n977);
	nor (gm_n3323, gm_n423, in_31, gm_n54, gm_n3322);
	or (gm_n3324, gm_n125, gm_n62, gm_n61, gm_n2274, gm_n314);
	or (gm_n3325, gm_n456, gm_n158, in_19, gm_n3324, gm_n514);
	nor (gm_n3326, gm_n583, in_31, gm_n54, gm_n3325, gm_n838);
	nor (gm_n3327, gm_n154, gm_n63, gm_n124, gm_n384, gm_n188);
	nand (gm_n3328, gm_n255, gm_n76, in_16, gm_n3327, gm_n270);
	nor (gm_n3329, gm_n248, gm_n83, in_24, gm_n3328, gm_n195);
	or (gm_n3330, gm_n670, gm_n62, in_11, gm_n621, gm_n398);
	or (gm_n3331, gm_n1225, in_23, in_19, gm_n3330, gm_n613);
	nor (gm_n3332, gm_n1112, gm_n55, in_27, gm_n3331, gm_n423);
	nand (gm_n3333, gm_n91, in_16, in_12, gm_n2012, gm_n340);
	or (gm_n3334, gm_n463, gm_n82, in_20, gm_n3333, gm_n411);
	nor (gm_n3335, gm_n185, gm_n85, in_28, gm_n3334);
	nand (gm_n3336, gm_n74, in_23, in_19, gm_n1106, gm_n77);
	nor (gm_n3337, gm_n977, in_31, gm_n54, gm_n3336, gm_n675);
	or (gm_n3338, gm_n3332, gm_n3329, gm_n3326, gm_n3337, gm_n3335);
	nand (gm_n3339, in_17, gm_n64, gm_n175, gm_n2723, gm_n2585);
	or (gm_n3340, gm_n1557, in_25, in_21, gm_n3339, gm_n1561);
	nor (gm_n3341, gm_n55, in_30, gm_n80, gm_n3340, gm_n3124);
	nor (gm_n3342, gm_n433, in_15, in_11, gm_n584, gm_n363);
	nand (gm_n3343, gm_n296, in_23, in_19, gm_n3342, gm_n1042);
	nor (gm_n3344, gm_n357, in_31, in_27, gm_n3343, gm_n977);
	nor (gm_n3345, gm_n599, in_12, gm_n124, gm_n298, gm_n971);
	and (gm_n3346, gm_n150, in_20, gm_n73, gm_n3345, gm_n270);
	and (gm_n3347, gm_n192, gm_n83, in_24, gm_n3346, gm_n215);
	and (gm_n3348, gm_n3347, gm_n101);
	or (gm_n3349, gm_n3348, gm_n3344, gm_n3341);
	nand (gm_n3350, gm_n150, gm_n63, gm_n124, gm_n1000, gm_n167);
	or (gm_n3351, gm_n187, gm_n76, gm_n73, gm_n3350, gm_n566);
	nor (gm_n3352, gm_n234, in_28, in_24, gm_n3351, gm_n248);
	and (gm_n3353, gm_n150, in_12, in_8, gm_n1946, gm_n256);
	nand (gm_n3354, gm_n107, gm_n76, in_16, gm_n3353, gm_n192);
	nor (gm_n3355, gm_n216, in_28, in_24, gm_n3354, gm_n226);
	and (gm_n3356, gm_n166, gm_n73, gm_n63, gm_n2514, gm_n228);
	nand (gm_n3357, gm_n255, in_24, in_20, gm_n3356, gm_n270);
	nor (gm_n3358, gm_n684, gm_n216, in_28, gm_n3357);
	or (gm_n3359, gm_n3358, gm_n3355, gm_n3352);
	or (gm_n3360, gm_n3338, gm_n3323, gm_n3320, gm_n3359, gm_n3349);
	nand (gm_n3361, gm_n299, gm_n62, in_11, gm_n394, gm_n698);
	or (gm_n3362, gm_n122, gm_n158, gm_n58, gm_n3361, gm_n317);
	nor (gm_n3363, gm_n423, gm_n55, gm_n54, gm_n3362, gm_n977);
	nand (gm_n3364, gm_n201, in_16, gm_n63, gm_n340, gm_n207);
	or (gm_n3365, gm_n520, gm_n82, gm_n76, gm_n3364, gm_n412);
	nor (gm_n3366, gm_n368, gm_n195, gm_n83, gm_n3365);
	nor (gm_n3367, gm_n93, gm_n63, gm_n124, gm_n288, gm_n168);
	and (gm_n3368, gm_n91, gm_n76, gm_n73, gm_n3367, gm_n235);
	and (gm_n3369, gm_n186, gm_n83, in_24, gm_n3368, gm_n263);
	and (gm_n3370, gm_n3369, gm_n196);
	or (gm_n3371, gm_n3370, gm_n3366, gm_n3363);
	nor (gm_n3372, gm_n374, in_16, gm_n63, gm_n1881, gm_n288);
	nand (gm_n3373, gm_n263, gm_n82, in_20, gm_n3372, gm_n477);
	nor (gm_n3374, gm_n224, gm_n185, gm_n83, gm_n3373);
	and (gm_n3375, in_7, gm_n115, gm_n70, gm_n361, in_8);
	and (gm_n3376, gm_n153, gm_n73, in_12, gm_n3375, gm_n446);
	and (gm_n3377, gm_n205, in_24, gm_n76, gm_n3376, gm_n477);
	and (gm_n3378, gm_n466, gm_n213, gm_n83, gm_n3377);
	nand (gm_n3379, gm_n199, in_12, in_8, gm_n1137, gm_n144);
	nor (gm_n3380, gm_n165, gm_n76, in_16, gm_n3379, gm_n236);
	nand (gm_n3381, gm_n186, gm_n83, gm_n82, gm_n3380, gm_n255);
	nor (gm_n3382, gm_n3381, gm_n479);
	or (gm_n3383, gm_n3382, gm_n3378, gm_n3374);
	or (gm_n3384, gm_n3360, gm_n3317, gm_n3314, gm_n3383, gm_n3371);
	nand (gm_n3385, gm_n167, gm_n73, in_12, gm_n1553, gm_n207);
	or (gm_n3386, gm_n566, in_24, gm_n76, gm_n3385, gm_n463);
	nor (gm_n3387, gm_n195, gm_n85, in_28, gm_n3386);
	nand (gm_n3388, gm_n392, gm_n62, in_11, gm_n2766, gm_n931);
	or (gm_n3389, gm_n1225, in_23, in_19, gm_n3388, gm_n1200);
	nor (gm_n3390, gm_n423, gm_n55, in_27, gm_n3389);
	nor (gm_n3391, gm_n393, gm_n58, in_15, gm_n2388, gm_n991);
	nand (gm_n3392, gm_n316, gm_n54, gm_n158, gm_n3391, gm_n459);
	nor (gm_n3393, gm_n3392, gm_n57, in_31);
	or (gm_n3394, gm_n3393, gm_n3390, gm_n3387);
	nor (gm_n3395, gm_n143, in_16, in_12, gm_n2070, gm_n599);
	nand (gm_n3396, gm_n107, gm_n82, in_20, gm_n3395, gm_n263);
	nor (gm_n3397, gm_n214, gm_n85, gm_n83, gm_n3396);
	and (gm_n3398, gm_n65, gm_n62, gm_n61, gm_n394, gm_n332);
	nand (gm_n3399, gm_n130, gm_n158, in_19, gm_n3398, gm_n1042);
	nor (gm_n3400, gm_n583, gm_n55, gm_n54, gm_n3399, gm_n675);
	and (gm_n3401, gm_n71, in_12, in_8, gm_n242, gm_n219);
	and (gm_n3402, gm_n446, in_20, gm_n73, gm_n3401, gm_n235);
	and (gm_n3403, gm_n139, gm_n83, in_24, gm_n3402, gm_n217);
	and (gm_n3404, gm_n3403, gm_n629);
	or (gm_n3405, gm_n3404, gm_n3400, gm_n3397);
	or (gm_n3406, gm_n3384, gm_n3311, gm_n3308, gm_n3405, gm_n3394);
	or (gm_n3407, gm_n796, gm_n62, in_11, gm_n1531, gm_n363);
	or (gm_n3408, gm_n1225, gm_n158, in_19, gm_n3407, gm_n422);
	nor (gm_n3409, gm_n423, in_31, gm_n54, gm_n3408);
	nand (gm_n3410, gm_n176, gm_n73, in_12, gm_n704, gm_n340);
	or (gm_n3411, gm_n566, in_24, in_20, gm_n3410, gm_n476);
	nor (gm_n3412, gm_n479, gm_n774, in_28, gm_n3411);
	nand (gm_n3413, gm_n176, in_20, in_16, gm_n1614, gm_n477);
	or (gm_n3414, gm_n89, in_28, in_24, gm_n3413, gm_n248);
	nor (gm_n3415, gm_n3414, gm_n195);
	or (gm_n3416, gm_n3415, gm_n3412, gm_n3409);
	nor (gm_n3417, gm_n92, in_15, in_8, gm_n1034, gm_n623);
	nand (gm_n3418, gm_n121, gm_n158, gm_n58, gm_n3417, gm_n173);
	nor (gm_n3419, gm_n1112, in_31, gm_n54, gm_n3418, gm_n612);
	and (gm_n3420, gm_n65, gm_n62, gm_n61, gm_n2581, gm_n995);
	nand (gm_n3421, gm_n296, gm_n158, in_19, gm_n3420, gm_n359);
	nor (gm_n3422, gm_n1200, gm_n55, gm_n54, gm_n3421, gm_n618);
	nor (gm_n3423, gm_n669, gm_n725, gm_n61, gm_n2141, gm_n447);
	and (gm_n3424, gm_n74, gm_n58, gm_n62, gm_n3423, gm_n316);
	and (gm_n3425, gm_n306, in_27, in_23, gm_n3424, gm_n657);
	and (gm_n3426, gm_n3425, in_31);
	or (gm_n3427, gm_n3426, gm_n3422, gm_n3419);
	or (gm_n3428, gm_n3406, gm_n3305, gm_n3301, gm_n3427, gm_n3416);
	nand (gm_n3429, gm_n1042, gm_n256, in_15, gm_n754, gm_n622);
	nor (gm_n3430, gm_n183, in_23, gm_n58, gm_n3429, gm_n335);
	nand (gm_n3431, gm_n438, gm_n55, gm_n54, gm_n3430);
	nor (gm_n3432, gm_n92, gm_n73, in_12, gm_n2543, gm_n177);
	and (gm_n3433, gm_n235, in_24, in_20, gm_n3432, gm_n263);
	nand (gm_n3434, gm_n213, gm_n84, in_28, gm_n3433);
	and (gm_n3435, gm_n153, gm_n63, gm_n124, gm_n402, gm_n515);
	nand (gm_n3436, gm_n1125, gm_n105, in_13, gm_n3435, gm_n2724);
	nor (gm_n3437, gm_n2209, in_25, in_21, gm_n3436, gm_n2182);
	nand (gm_n3438, gm_n55, gm_n100, gm_n80, gm_n3437);
	nand (gm_n3439, gm_n3438, gm_n3434, gm_n3431);
	or (gm_n3440, gm_n599, gm_n73, in_12, gm_n3104, gm_n177);
	nor (gm_n3441, gm_n197, in_24, in_20, gm_n3440, gm_n630);
	nand (gm_n3442, gm_n186, gm_n81, in_28, gm_n3441);
	nand (gm_n3443, gm_n166, in_20, gm_n73, gm_n1191, gm_n235);
	nor (gm_n3444, gm_n630, in_28, gm_n82, gm_n3443, gm_n368);
	nand (gm_n3445, gm_n3444, gm_n137);
	nand (gm_n3446, gm_n91, in_16, gm_n63, gm_n589, gm_n199);
	nor (gm_n3447, gm_n165, gm_n82, gm_n76, gm_n3446, gm_n520);
	nand (gm_n3448, gm_n466, gm_n196, gm_n83, gm_n3447);
	nand (gm_n3449, gm_n3448, gm_n3445, gm_n3442);
	or (gm_n3450, gm_n3428, gm_n3298, gm_n3295, gm_n3449, gm_n3439);
	nor (gm_n3451, gm_n796, in_15, gm_n61, gm_n2795, gm_n991);
	and (gm_n3452, gm_n134, gm_n158, gm_n58, gm_n3451, gm_n334);
	and (gm_n3453, gm_n438, in_31, in_27, gm_n3452);
	and (gm_n3454, gm_n65, gm_n62, gm_n61, gm_n1710, gm_n995);
	and (gm_n3455, gm_n121, in_23, in_19, gm_n3454, gm_n358);
	and (gm_n3456, gm_n337, gm_n55, in_27, gm_n3455, gm_n459);
	nor (gm_n3457, gm_n553, in_12, in_8, gm_n1034, gm_n288);
	nand (gm_n3458, gm_n235, in_20, gm_n73, gm_n3457, gm_n255);
	nor (gm_n3459, gm_n185, in_28, in_24, gm_n3458, gm_n262);
	nor (gm_n3460, gm_n3459, gm_n3456, gm_n3453);
	not (gm_n3461, gm_n3460);
	and (gm_n3462, gm_n446, in_16, in_12, gm_n2205, gm_n228);
	and (gm_n3463, gm_n227, in_24, in_20, gm_n3462, gm_n235);
	and (gm_n3464, gm_n367, gm_n213, gm_n83, gm_n3463);
	or (gm_n3465, gm_n3450, gm_n3292, gm_n3289, gm_n3464, gm_n3461);
	nand (gm_n3466, gm_n3465, gm_n3288);
	nand (new_out1, gm_n3466, gm_n3109);
	and (new_out2, gm_n3288, gm_n2930);
	and (new_out3, gm_n3465, gm_n3108);
	nand (new_out4, gm_n3465, gm_n2930);
	nor (new_out5, gm_n3288, gm_n3108);
endmodule

module top ( g0 , g1 , g2 , g3 , g4 , g5 , g6 , g7 , g8 , g9 , g10 , g11 , g12 , g13 , g14 , g15 , g16 , g17 , g18 , g19 , g20 , g21 , g22 , g23 , g24 , g25 , g26 , g27 , g28 , g29 , g30 , g31 , g32 , g33 , g34 , g35 , g36 , g37 , g38 , g39 , g40 , g41 , g42 , g43 , g44 , g45 , g46 , g47 , g48 , g49 , g50 , g51 , g52 , g53 , g54 , g55 , g56 , g57 , g58 , g59 , g60 , g61 , g62 , g63 , g64 , g65 , g66 , g67 , g68 , g69 , g70 , g71 , g72 , g73 , g74 , g75 , g76 , g77 , g78 , g79 , g80 , g81 , g82 , g83 , g84 , g85 , g86 , g87 , g88 , g89 , g90 , g91 , g92 , g93 , g94 , g95 , g96 , g97 , g98 , g99 , g100 , g101 , g102 , g103 , g104 , g105 , g106 , g107 , g108 , g109 , g110 , g111 , g112 , g113 , g114 , g115 , g116 , g117 , g118 , g119 , g120 , g121 , g122 , g123 , g124 , g125 , g126 , g127 , g128 , g129 , g130 , g131 , g132 , g133 , g134 , g135 , g136 , g137 , g138 , g139 , g140 , g141 , g142 , g143 , g144 , g145 , g146 , g147 , g148 , g149 , g150 , g151 , g152 , g153 , g154 , g155 , g156 , g157 , g158 , g159 , g160 , g161 , g162 , g163 , g164 , g165 , g166 , g167 , g168 , g169 , g170 , g171 , g172 , g173 , g174 , g175 , g176 , g177 , g178 , g179 , g180 , g181 , g182 , g183 , g184 , g185 , g186 , g187 , g188 , g189 , g190 , g191 , g192 , g193 , g194 , g195 , g196 , g197 , g198 , g199 , g200 , g201 , g202 , g203 , g204 , g205 , g206 , g207 , g208 , g209 , g210 , g211 , g212 , g213 , g214 , g215 , g216 , g217 , g218 , g219 , g220 , g221 , g222 , g223 , g224 , g225 , g226 , g227 , g228 , g229 , g230 , g231 , g232 , g233 , g234 , g235 , g236 , g237 , g238 , g239 , g240 , g241 , g242 , g243 , g244 , g245 , g246 , g247 , g248 , g249 , g250 , g251 , g252 , g253 , g254 , g255 , g256 , g257 , g258 , g259 , g260 , g261 , g262 , g263 , g264 , g265 , g266 , g267 , g268 , g269 , g270 , g271 , g272 , g273 , g274 , g275 , g276 , g277 , g278 , g279 , g280 , g281 , g282 , g283 , g284 , g285 , g286 , g287 , g288 , g289 , g290 , g291 , g292 , g293 , g294 , g295 , g296 , g297 , g298 , g299 , g300 , g301 , g302 , g303 , g304 , g305 , g306 , g307 , g308 , g309 , g310 , g311 , g312 , g313 , g314 , g315 , g316 , g317 , g318 , g319 , g320 , g321 , g322 , g323 , g324 , g325 , g326 , g327 , g328 , g329 , g330 , g331 , g332 , g333 , g334 , g335 , g336 , g337 , g338 , g339 , g340 , g341 , g342 , g343 , g344 , g345 , g346 , g347 , g348 , g349 , g350 , g351 , g352 , g353 , g354 , g355 , g356 , g357 , g358 , g359 , g360 , g361 , g362 , g363 , g364 , g365 , g366 , g367 , g368 , g369 , g370 , g371 , g372 , g373 , g374 , g375 , g376 , g377 , g378 , g379 , g380 , g381 , g382 , g383 , g384 , g385 , g386 , g387 , g388 , g389 , g390 , g391 , g392 , g393 , g394 , g395 , g396 , g397 , g398 , g399 , g400 , g401 , g402 , g403 , g404 , g405 , g406 , g407 , g408 , g409 , g410 , new_out1, new_out2, new_out3, new_out4, new_out5 );
	input g0, g1, g2, g3, g4, g5, g6, g7, g8, g9, g10, g11, g12, g13, g14, g15, g16, g17, g18, g19, g20, g21, g22, g23, g24, g25, g26, g27, g28, g29, g30, g31, g32, g33, g34, g35, g36, g37, g38, g39, g40, g41, g42, g43, g44, g45, g46, g47, g48, g49, g50, g51, g52, g53, g54, g55, g56, g57, g58, g59, g60, g61, g62, g63, g64, g65, g66, g67, g68, g69, g70, g71, g72, g73, g74, g75, g76, g77, g78, g79, g80, g81, g82, g83, g84, g85, g86, g87, g88, g89, g90, g91, g92, g93, g94, g95, g96, g97, g98, g99, g100, g101, g102, g103, g104, g105, g106, g107, g108, g109, g110, g111, g112, g113, g114, g115, g116, g117, g118, g119, g120, g121, g122, g123, g124, g125, g126, g127, g128, g129, g130, g131, g132, g133, g134, g135, g136, g137, g138, g139, g140, g141, g142, g143, g144, g145, g146, g147, g148, g149, g150, g151, g152, g153, g154, g155, g156, g157, g158, g159, g160, g161, g162, g163, g164, g165, g166, g167, g168, g169, g170, g171, g172, g173, g174, g175, g176, g177, g178, g179, g180, g181, g182, g183, g184, g185, g186, g187, g188, g189, g190, g191, g192, g193, g194, g195, g196, g197, g198, g199, g200, g201, g202, g203, g204, g205, g206, g207, g208, g209, g210, g211, g212, g213, g214, g215, g216, g217, g218, g219, g220, g221, g222, g223, g224, g225, g226, g227, g228, g229, g230, g231, g232, g233, g234, g235, g236, g237, g238, g239, g240, g241, g242, g243, g244, g245, g246, g247, g248, g249, g250, g251, g252, g253, g254, g255, g256, g257, g258, g259, g260, g261, g262, g263, g264, g265, g266, g267, g268, g269, g270, g271, g272, g273, g274, g275, g276, g277, g278, g279, g280, g281, g282, g283, g284, g285, g286, g287, g288, g289, g290, g291, g292, g293, g294, g295, g296, g297, g298, g299, g300, g301, g302, g303, g304, g305, g306, g307, g308, g309, g310, g311, g312, g313, g314, g315, g316, g317, g318, g319, g320, g321, g322, g323, g324, g325, g326, g327, g328, g329, g330, g331, g332, g333, g334, g335, g336, g337, g338, g339, g340, g341, g342, g343, g344, g345, g346, g347, g348, g349, g350, g351, g352, g353, g354, g355, g356, g357, g358, g359, g360, g361, g362, g363, g364, g365, g366, g367, g368, g369, g370, g371, g372, g373, g374, g375, g376, g377, g378, g379, g380, g381, g382, g383, g384, g385, g386, g387, g388, g389, g390, g391, g392, g393, g394, g395, g396, g397, g398, g399, g400, g401, g402, g403, g404, g405, g406, g407, g408, g409, g410;
	output new_out1, new_out2, new_out3, new_out4, new_out5;
	wire gm_n421, gm_n422, gm_n423, gm_n424, gm_n426, gm_n427, gm_n428, gm_n430, gm_n431, gm_n432, gm_n433, gm_n435, gm_n436, gm_n437, gm_n439;
	wire t_3, t_1, t_0, t_2;
	and (gm_n421, g401, g370);
	not (gm_n422, g370);
	and (gm_n423, g400, gm_n422);
	or (gm_n424, gm_n423, gm_n421);
	and (new_out2, gm_n424, t_0);
	and (gm_n426, g404, g370);
	and (gm_n427, g403, gm_n422);
	or (gm_n428, gm_n427, gm_n426);
	and (new_out3, gm_n428, t_1);
	or (gm_n430, new_out3, new_out2);
	and (gm_n431, g370, g5);
	and (gm_n432, g407, gm_n422);
	or (gm_n433, gm_n432, gm_n431);
	and (new_out4, gm_n433, t_2);
	and (gm_n435, g370, g4);
	and (gm_n436, g410, gm_n422);
	or (gm_n437, gm_n436, gm_n435);
	and (new_out5, gm_n437, t_3);
	or (gm_n439, new_out5, new_out4);
	nand (new_out1, gm_n439, gm_n430);
endmodule
